library IEEE;

use IEEE.std_logic_1164.all;
-- use ieee.numeric_std.all;

package 
   CONV_PACK 
   is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type UNSIGNED is array (INTEGER range <>) of std_logic;
   
   -- Declarations for conversion functions.
   function BIT_to_std_logic(arg : in BIT) return std_logic;

end 
   CONV_PACK;

package body 
   CONV_PACK 
   is
   
   -- enum type to std_logic function
   function BIT_to_std_logic(arg : in BIT) return std_logic is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when '0' => return '0';
         when '1' => return '1';
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return '0';
      end case;
   end;

end 
   CONV_PACK;

library IEEE;

use IEEE.std_logic_1164.all;

use 
   work.CONV_PACK.all;

entity 
   top_g_hub_mux3_g_clock_freq200000000_g_color_depth8_g_num_row4_g_num_col8_g_addr_width5_g_u_row2_g_u_col3 
   is

   port( clk : in std_logic;  reset : in bit;  top_data : in bit_vector 
         (23 downto 0);  top_dv_i, top_u_l : in bit;  top_ack : out 
         bit;  hub_mux_o : out bit_vector (2 downto 0);  hub_clk_o, 
         hub_latch_o, hub_blank_o, hub_g0_o, hub_b0_o, hub_r0_o : out bit
         );

end 
   top_g_hub_mux3_g_clock_freq200000000_g_color_depth8_g_num_row4_g_num_col8_g_addr_width5_g_u_row2_g_u_col3;

architecture SYN_rtl of 
   top_g_hub_mux3_g_clock_freq200000000_g_color_depth8_g_num_row4_g_num_col8_g_addr_width5_g_u_row2_g_u_col3 
   is

   component inv
      port( inb : in bit;  outb : out bit);
   end component;
   
   component nand3
      port( a, b, c : in bit;  outb : out bit);
   end component;
   
   component nand2
      port( a, b : in bit;  outb : out bit);
   end component;
   
   component oai12
      port( b, c, a : in bit;  outb : out bit);
   end component;
   
   component nor3
      port( a, b, c : in bit;  outb : out bit);
   end component;
   
   component nor2
      port( a, b : in bit;  outb : out bit);
   end component;
   
   component aoi12
      port( b, c, a : in bit;  outb : out bit);
   end component;
   
   component oai22
      port( a, b, c, d : in bit;  outb : out bit);
   end component;
   
   component nand4
      port( a, b, c, d : in bit;  outb : out bit);
   end component;
   
   component aoi22
      port( a, b, c, d : in bit;  outb : out bit);
   end component;
   
   component xor2
      port( a, b : in bit;  outb : out bit);
   end component;
   
   component dff
      port( gclk: in std_logic; d, rnot: in bit;  q : out bit);
   end component;
   
   signal reset_port, top_ack_port, hub_mux_o_2_port, hub_mux_o_1_port, 
      hub_mux_o_0_port, hub_clk_o_port, hub_latch_o_port, hub_blank_o_port, 
      hub_g0_o_port, hub_b0_o_port, hub_r0_o_port, mem_sipo_r0_7_port, 
      mem_sipo_r0_6_port, mem_sipo_r0_5_port, mem_sipo_r0_4_port, 
      mem_sipo_r0_3_port, mem_sipo_r0_2_port, mem_sipo_r0_1_port, 
      mem_sipo_r0_0_port, mem_sipo_g0_7_port, mem_sipo_g0_6_port, 
      mem_sipo_g0_5_port, mem_sipo_g0_4_port, mem_sipo_g0_3_port, 
      mem_sipo_g0_2_port, mem_sipo_g0_1_port, mem_sipo_g0_0_port, 
      mem_sipo_b0_7_port, mem_sipo_b0_6_port, mem_sipo_b0_5_port, 
      mem_sipo_b0_4_port, mem_sipo_b0_3_port, mem_sipo_b0_2_port, 
      mem_sipo_b0_1_port, mem_sipo_b0_0_port, mem_out_r0_7_port, 
      mem_out_r0_6_port, mem_out_r0_5_port, mem_out_r0_4_port, 
      mem_out_r0_3_port, mem_out_r0_2_port, mem_out_r0_1_port, 
      mem_out_r0_0_port, mem_out_g0_7_port, mem_out_g0_6_port, 
      mem_out_g0_5_port, mem_out_g0_4_port, mem_out_g0_3_port, 
      mem_out_g0_2_port, mem_out_g0_1_port, mem_out_g0_0_port, 
      mem_out_b0_7_port, mem_out_b0_6_port, mem_out_b0_5_port, 
      mem_out_b0_4_port, mem_out_b0_3_port, mem_out_b0_2_port, 
      mem_out_b0_1_port, mem_out_b0_0_port, addr_i_4_port, addr_i_3_port, 
      addr_i_2_port, addr_i_1_port, addr_i_0_port, reg_hub_f, hub_reg_f, 
      mem_reg_f, mem_hub_f, registers_n296, registers_n295, registers_n294, 
      registers_n293, registers_n292, registers_n291, registers_n290, 
      registers_n289, registers_n288, registers_n287, registers_n286, 
      registers_n285, registers_n284, registers_n283, registers_n282, 
      registers_n281, registers_n280, registers_n279, registers_n278, 
      registers_n277, registers_n276, registers_n275, registers_n274, 
      registers_n273, registers_n272, registers_n271, registers_n270, 
      registers_n269, registers_n268, registers_n267, registers_n266, 
      registers_n265, registers_n264, registers_n263, registers_n262, 
      registers_n261, registers_n260, registers_n259, registers_n258, 
      registers_n257, registers_n256, registers_n255, registers_n254, 
      registers_n253, registers_n252, registers_n251, registers_n250, 
      registers_n249, registers_n248, registers_n247, registers_n246, 
      registers_n245, registers_n244, registers_n243, registers_n242, 
      registers_n241, registers_n240, registers_n239, registers_n238, 
      registers_n237, registers_n236, registers_n235, registers_n234, 
      registers_n233, registers_n232, registers_n84, registers_n83, 
      registers_n82, registers_n81, registers_n80, registers_n79, registers_n78
      , registers_n77, registers_n76, registers_n75, registers_n74, 
      registers_n73, registers_n72, registers_n71, registers_n70, registers_n69
      , registers_n68, registers_n67, registers_n66, registers_n65, 
      registers_n64, registers_n63, registers_n62, registers_n61, registers_n60
      , registers_n59, registers_n58, registers_n57, registers_n56, 
      registers_n55, registers_n54, registers_n53, registers_n52, registers_n51
      , registers_n50, registers_n49, registers_n48, registers_n47, 
      registers_n46, registers_n45, registers_n44, registers_n43, registers_n42
      , registers_n41, registers_n40, registers_n39, registers_n38, 
      registers_n37, registers_n36, registers_n35, registers_n34, registers_n33
      , registers_n32, registers_n31, registers_n30, registers_n29, 
      registers_n28, registers_n27, registers_n26, registers_n25, registers_n24
      , registers_n23, registers_n22, registers_n21, registers_n20, 
      registers_n19, registers_s_delay_0_port, registers_s_delay_1_port, 
      registers_s_mem_sipo_b0_0_port, registers_s_mem_sipo_b0_1_port, 
      registers_s_mem_sipo_b0_2_port, registers_s_mem_sipo_b0_3_port, 
      registers_s_mem_sipo_b0_4_port, registers_s_mem_sipo_b0_5_port, 
      registers_s_mem_sipo_b0_6_port, registers_s_mem_sipo_b0_7_port, 
      registers_s_mem_sipo_g0_0_port, registers_s_mem_sipo_g0_1_port, 
      registers_s_mem_sipo_g0_2_port, registers_s_mem_sipo_g0_3_port, 
      registers_s_mem_sipo_g0_4_port, registers_s_mem_sipo_g0_5_port, 
      registers_s_mem_sipo_g0_6_port, registers_s_mem_sipo_g0_7_port, 
      registers_s_mem_sipo_r0_0_port, registers_s_mem_sipo_r0_1_port, 
      registers_s_mem_sipo_r0_2_port, registers_s_mem_sipo_r0_3_port, 
      registers_s_mem_sipo_r0_4_port, registers_s_mem_sipo_r0_5_port, 
      registers_s_mem_sipo_r0_6_port, registers_s_mem_sipo_r0_7_port, 
      registers_reg_col_inc_0_port, registers_reg_col_inc_1_port, 
      registers_reg_col_inc_2_port, registers_reg_cd_0_port, 
      registers_reg_cd_1_port, registers_reg_cd_2_port, 
      registers_reg_row_0_port, registers_reg_row_1_port, 
      registers_mem_to_reg_0_port, registers_mem_to_reg_1_port, 
      load_n_store_n275, load_n_store_n274, load_n_store_n273, 
      load_n_store_n272, load_n_store_n271, load_n_store_n270, 
      load_n_store_n269, load_n_store_n268, load_n_store_n267, 
      load_n_store_n266, load_n_store_n265, load_n_store_n264, 
      load_n_store_n263, load_n_store_n262, load_n_store_n261, 
      load_n_store_n260, load_n_store_n259, load_n_store_n76, load_n_store_n75,
      load_n_store_n74, load_n_store_n73, load_n_store_n72, load_n_store_n71, 
      load_n_store_n70, load_n_store_n69, load_n_store_n68, load_n_store_n67, 
      load_n_store_n66, load_n_store_n65, load_n_store_n64, load_n_store_n63, 
      load_n_store_n62, load_n_store_n61, load_n_store_n60, load_n_store_n59, 
      load_n_store_n58, load_n_store_n57, load_n_store_n56, load_n_store_n55, 
      load_n_store_n54, load_n_store_n53, load_n_store_n52, load_n_store_n51, 
      load_n_store_n50, load_n_store_n49, load_n_store_n48, load_n_store_n47, 
      load_n_store_n46, load_n_store_n45, load_n_store_n44, load_n_store_n43, 
      load_n_store_n42, load_n_store_n41, load_n_store_n40, load_n_store_n39, 
      load_n_store_n38, load_n_store_n37, load_n_store_n36, load_n_store_n35, 
      load_n_store_n34, load_n_store_n33, load_n_store_n32, load_n_store_n31, 
      load_n_store_n30, load_n_store_n29, load_n_store_n28, load_n_store_n27, 
      load_n_store_n26, load_n_store_n25, load_n_store_n24, load_n_store_n23, 
      load_n_store_n22, load_n_store_n21, load_n_store_n20, load_n_store_n19, 
      load_n_store_n18, load_n_store_n17, load_n_store_n16, load_n_store_n15, 
      load_n_store_n14, load_n_store_n13, load_n_store_n12, 
      load_n_store_mem_timer_0_port, load_n_store_mem_timer_1_port, 
      load_n_store_mem_timer_2_port, load_n_store_mem_timer_3_port, 
      load_n_store_mem_timer_4_port, load_n_store_mem_full, 
      load_n_store_simple_mem_sm_0_port, load_n_store_simple_mem_sm_1_port, 
      load_n_store_lazy_in_2_0_port, load_n_store_lazy_in_2_1_port, 
      load_n_store_lazy_in_2_2_port, load_n_store_lazy_in_2_3_port, 
      load_n_store_lazy_in_2_4_port, load_n_store_lazy_in_2_5_port, 
      load_n_store_lazy_in_2_6_port, load_n_store_lazy_in_2_7_port, 
      load_n_store_lazy_in_1_0_port, load_n_store_lazy_in_1_1_port, 
      load_n_store_lazy_in_1_2_port, load_n_store_lazy_in_1_3_port, 
      load_n_store_lazy_in_1_4_port, load_n_store_lazy_in_1_5_port, 
      load_n_store_lazy_in_1_6_port, load_n_store_lazy_in_1_7_port, 
      load_n_store_lazy_in_0_0_port, load_n_store_lazy_in_0_1_port, 
      load_n_store_lazy_in_0_2_port, load_n_store_lazy_in_0_3_port, 
      load_n_store_lazy_in_0_4_port, load_n_store_lazy_in_0_5_port, 
      load_n_store_lazy_in_0_6_port, load_n_store_lazy_in_0_7_port, 
      load_n_store_lazy_out_2_0_port, load_n_store_lazy_out_2_1_port, 
      load_n_store_lazy_out_2_2_port, load_n_store_lazy_out_2_3_port, 
      load_n_store_lazy_out_2_4_port, load_n_store_lazy_out_2_5_port, 
      load_n_store_lazy_out_2_6_port, load_n_store_lazy_out_2_7_port, 
      load_n_store_lazy_out_1_0_port, load_n_store_lazy_out_1_1_port, 
      load_n_store_lazy_out_1_2_port, load_n_store_lazy_out_1_3_port, 
      load_n_store_lazy_out_1_4_port, load_n_store_lazy_out_1_5_port, 
      load_n_store_lazy_out_1_6_port, load_n_store_lazy_out_1_7_port, 
      load_n_store_lazy_out_0_0_port, load_n_store_lazy_out_0_1_port, 
      load_n_store_lazy_out_0_2_port, load_n_store_lazy_out_0_3_port, 
      load_n_store_lazy_out_0_4_port, load_n_store_lazy_out_0_5_port, 
      load_n_store_lazy_out_0_6_port, load_n_store_lazy_out_0_7_port, 
      load_n_store_s_addr_0_port, load_n_store_s_addr_1_port, 
      load_n_store_s_addr_2_port, load_n_store_s_addr_3_port, 
      load_n_store_s_addr_4_port, load_n_store_we_i, display_out_n535, 
      display_out_n534, display_out_n533, display_out_n532, display_out_n531, 
      display_out_n530, display_out_n529, display_out_n528, display_out_n527, 
      display_out_n526, display_out_n525, display_out_n524, display_out_n523, 
      display_out_n522, display_out_n521, display_out_n520, display_out_n519, 
      display_out_n518, display_out_n517, display_out_n516, display_out_n515, 
      display_out_n514, display_out_n513, display_out_n512, display_out_n511, 
      display_out_n510, display_out_n509, display_out_n508, display_out_n507, 
      display_out_n506, display_out_n505, display_out_n504, display_out_n503, 
      display_out_n502, display_out_n501, display_out_n500, display_out_n499, 
      display_out_n498, display_out_n497, display_out_n496, display_out_n495, 
      display_out_n494, display_out_n493, display_out_n492, display_out_n491, 
      display_out_n490, display_out_n489, display_out_n488, display_out_n487, 
      display_out_n486, display_out_n485, display_out_n484, display_out_n483, 
      display_out_n482, display_out_n481, display_out_n480, display_out_n479, 
      display_out_n478, display_out_n477, display_out_n476, display_out_n475, 
      display_out_n474, display_out_n151, display_out_n150, display_out_n149, 
      display_out_n148, display_out_n147, display_out_n146, display_out_n145, 
      display_out_n144, display_out_n143, display_out_n142, display_out_n141, 
      display_out_n140, display_out_n139, display_out_n138, display_out_n137, 
      display_out_n136, display_out_n135, display_out_n134, display_out_n133, 
      display_out_n132, display_out_n131, display_out_n130, display_out_n129, 
      display_out_n128, display_out_n127, display_out_n126, display_out_n125, 
      display_out_n124, display_out_n123, display_out_n122, display_out_n121, 
      display_out_n120, display_out_n119, display_out_n118, display_out_n117, 
      display_out_n116, display_out_n115, display_out_n114, display_out_n113, 
      display_out_n112, display_out_n111, display_out_n110, display_out_n109, 
      display_out_n108, display_out_n107, display_out_n106, display_out_n105, 
      display_out_n104, display_out_n103, display_out_n102, display_out_n101, 
      display_out_n100, display_out_n99, display_out_n98, display_out_n97, 
      display_out_n96, display_out_n95, display_out_n94, display_out_n93, 
      display_out_n92, display_out_n91, display_out_n90, display_out_n89, 
      display_out_n88, display_out_n87, display_out_n86, display_out_n85, 
      display_out_n84, display_out_n83, display_out_n82, display_out_n81, 
      display_out_n80, display_out_n79, display_out_n78, display_out_n77, 
      display_out_n76, display_out_n75, display_out_n74, display_out_n73, 
      display_out_n72, display_out_n71, display_out_n70, display_out_n69, 
      display_out_n68, display_out_hub_piso_b0_0_port, 
      display_out_hub_piso_b0_1_port, display_out_hub_piso_b0_2_port, 
      display_out_hub_piso_b0_3_port, display_out_hub_piso_b0_4_port, 
      display_out_hub_piso_b0_5_port, display_out_hub_piso_b0_6_port, 
      display_out_hub_piso_b0_7_port, display_out_hub_piso_g0_0_port, 
      display_out_hub_piso_g0_1_port, display_out_hub_piso_g0_2_port, 
      display_out_hub_piso_g0_3_port, display_out_hub_piso_g0_4_port, 
      display_out_hub_piso_g0_5_port, display_out_hub_piso_g0_6_port, 
      display_out_hub_piso_g0_7_port, display_out_hub_piso_r0_0_port, 
      display_out_hub_piso_r0_1_port, display_out_hub_piso_r0_2_port, 
      display_out_hub_piso_r0_3_port, display_out_hub_piso_r0_4_port, 
      display_out_hub_piso_r0_5_port, display_out_hub_piso_r0_6_port, 
      display_out_hub_piso_r0_7_port, display_out_clk_timer_0_port, 
      display_out_clk_timer_1_port, display_out_clk_timer_2_port, 
      display_out_clk_timer_3_port, display_out_clk_timer_4_port, 
      display_out_clk_timer_5_port, display_out_clk_timer_6_port, 
      display_out_disp_timer_0_port, display_out_disp_timer_1_port, 
      display_out_disp_timer_2_port, display_out_disp_timer_3_port, 
      display_out_disp_timer_4_port, display_out_disp_timer_5_port, 
      display_out_disp_timer_6_port, display_out_disp_timer_7_port, 
      display_out_disp_timer_8_port, display_out_disp_timer_9_port, 
      display_out_disp_timer_10_port, display_out_disp_timer_11_port, 
      display_out_disp_timer_12_port, display_out_disp_timer_13_port, 
      display_out_disp_timer_14_port, display_out_disp_timer_15_port, 
      display_out_disp_timer_16_port, display_out_disp_timer_17_port, 
      display_out_disp_timer_18_port, display_out_disp_timer_19_port, 
      display_out_disp_timer_20_port, display_out_disp_timer_21_port, 
      display_out_disp_timer_22_port, display_out_disp_timer_23_port, 
      display_out_disp_timer_24_port, display_out_disp_timer_25_port, 
      display_out_disp_timer_26_port, display_out_disp_timer_27_port, 
      display_out_disp_timer_28_port, display_out_disp_timer_29_port, 
      display_out_disp_timer_30_port, display_out_disp_timer_31_port, 
      display_out_h_col_0_port, display_out_h_col_1_port, 
      display_out_h_col_2_port, display_out_h_row_0_port, 
      display_out_h_row_1_port, display_out_bcd_time_0_port, 
      display_out_bcd_time_1_port, display_out_bcd_time_2_port, 
      display_out_hub_out_sm_0_port, display_out_hub_out_sm_1_port, 
      display_out_hub_out_sm_2_port, load_n_store_RGB_Array_0_n1162, 
      load_n_store_RGB_Array_0_n1161, load_n_store_RGB_Array_0_n1160, 
      load_n_store_RGB_Array_0_n1159, load_n_store_RGB_Array_0_n1158, 
      load_n_store_RGB_Array_0_n1157, load_n_store_RGB_Array_0_n1156, 
      load_n_store_RGB_Array_0_n1155, load_n_store_RGB_Array_0_n1154, 
      load_n_store_RGB_Array_0_n1153, load_n_store_RGB_Array_0_n1152, 
      load_n_store_RGB_Array_0_n1151, load_n_store_RGB_Array_0_n1150, 
      load_n_store_RGB_Array_0_n1149, load_n_store_RGB_Array_0_n1148, 
      load_n_store_RGB_Array_0_n1147, load_n_store_RGB_Array_0_n1146, 
      load_n_store_RGB_Array_0_n1145, load_n_store_RGB_Array_0_n1144, 
      load_n_store_RGB_Array_0_n1143, load_n_store_RGB_Array_0_n1142, 
      load_n_store_RGB_Array_0_n1141, load_n_store_RGB_Array_0_n1140, 
      load_n_store_RGB_Array_0_n1139, load_n_store_RGB_Array_0_n1138, 
      load_n_store_RGB_Array_0_n1137, load_n_store_RGB_Array_0_n1136, 
      load_n_store_RGB_Array_0_n1135, load_n_store_RGB_Array_0_n1134, 
      load_n_store_RGB_Array_0_n1133, load_n_store_RGB_Array_0_n1132, 
      load_n_store_RGB_Array_0_n1131, load_n_store_RGB_Array_0_n1130, 
      load_n_store_RGB_Array_0_n1129, load_n_store_RGB_Array_0_n1128, 
      load_n_store_RGB_Array_0_n1127, load_n_store_RGB_Array_0_n1126, 
      load_n_store_RGB_Array_0_n1125, load_n_store_RGB_Array_0_n1124, 
      load_n_store_RGB_Array_0_n1123, load_n_store_RGB_Array_0_n1122, 
      load_n_store_RGB_Array_0_n1121, load_n_store_RGB_Array_0_n1120, 
      load_n_store_RGB_Array_0_n1119, load_n_store_RGB_Array_0_n1118, 
      load_n_store_RGB_Array_0_n1117, load_n_store_RGB_Array_0_n1116, 
      load_n_store_RGB_Array_0_n1115, load_n_store_RGB_Array_0_n1114, 
      load_n_store_RGB_Array_0_n1113, load_n_store_RGB_Array_0_n1112, 
      load_n_store_RGB_Array_0_n1111, load_n_store_RGB_Array_0_n1110, 
      load_n_store_RGB_Array_0_n1109, load_n_store_RGB_Array_0_n1108, 
      load_n_store_RGB_Array_0_n1107, load_n_store_RGB_Array_0_n1106, 
      load_n_store_RGB_Array_0_n1105, load_n_store_RGB_Array_0_n1104, 
      load_n_store_RGB_Array_0_n1103, load_n_store_RGB_Array_0_n1102, 
      load_n_store_RGB_Array_0_n1101, load_n_store_RGB_Array_0_n1100, 
      load_n_store_RGB_Array_0_n1099, load_n_store_RGB_Array_0_n1098, 
      load_n_store_RGB_Array_0_n1097, load_n_store_RGB_Array_0_n1096, 
      load_n_store_RGB_Array_0_n1095, load_n_store_RGB_Array_0_n1094, 
      load_n_store_RGB_Array_0_n1093, load_n_store_RGB_Array_0_n1092, 
      load_n_store_RGB_Array_0_n1091, load_n_store_RGB_Array_0_n1090, 
      load_n_store_RGB_Array_0_n1089, load_n_store_RGB_Array_0_n1088, 
      load_n_store_RGB_Array_0_n1087, load_n_store_RGB_Array_0_n1086, 
      load_n_store_RGB_Array_0_n1085, load_n_store_RGB_Array_0_n1084, 
      load_n_store_RGB_Array_0_n1083, load_n_store_RGB_Array_0_n1082, 
      load_n_store_RGB_Array_0_n1081, load_n_store_RGB_Array_0_n1080, 
      load_n_store_RGB_Array_0_n1079, load_n_store_RGB_Array_0_n1078, 
      load_n_store_RGB_Array_0_n1077, load_n_store_RGB_Array_0_n1076, 
      load_n_store_RGB_Array_0_n1075, load_n_store_RGB_Array_0_n1074, 
      load_n_store_RGB_Array_0_n1073, load_n_store_RGB_Array_0_n1072, 
      load_n_store_RGB_Array_0_n1071, load_n_store_RGB_Array_0_n1070, 
      load_n_store_RGB_Array_0_n1069, load_n_store_RGB_Array_0_n1068, 
      load_n_store_RGB_Array_0_n1067, load_n_store_RGB_Array_0_n1066, 
      load_n_store_RGB_Array_0_n1065, load_n_store_RGB_Array_0_n1064, 
      load_n_store_RGB_Array_0_n1063, load_n_store_RGB_Array_0_n1062, 
      load_n_store_RGB_Array_0_n1061, load_n_store_RGB_Array_0_n1060, 
      load_n_store_RGB_Array_0_n1059, load_n_store_RGB_Array_0_n1058, 
      load_n_store_RGB_Array_0_n1057, load_n_store_RGB_Array_0_n1056, 
      load_n_store_RGB_Array_0_n1055, load_n_store_RGB_Array_0_n1054, 
      load_n_store_RGB_Array_0_n1053, load_n_store_RGB_Array_0_n1052, 
      load_n_store_RGB_Array_0_n1051, load_n_store_RGB_Array_0_n1050, 
      load_n_store_RGB_Array_0_n1049, load_n_store_RGB_Array_0_n1048, 
      load_n_store_RGB_Array_0_n1047, load_n_store_RGB_Array_0_n1046, 
      load_n_store_RGB_Array_0_n1045, load_n_store_RGB_Array_0_n1044, 
      load_n_store_RGB_Array_0_n1043, load_n_store_RGB_Array_0_n1042, 
      load_n_store_RGB_Array_0_n1041, load_n_store_RGB_Array_0_n1040, 
      load_n_store_RGB_Array_0_n1039, load_n_store_RGB_Array_0_n1038, 
      load_n_store_RGB_Array_0_n1037, load_n_store_RGB_Array_0_n1036, 
      load_n_store_RGB_Array_0_n1035, load_n_store_RGB_Array_0_n1034, 
      load_n_store_RGB_Array_0_n1033, load_n_store_RGB_Array_0_n1032, 
      load_n_store_RGB_Array_0_n1031, load_n_store_RGB_Array_0_n1030, 
      load_n_store_RGB_Array_0_n1029, load_n_store_RGB_Array_0_n1028, 
      load_n_store_RGB_Array_0_n1027, load_n_store_RGB_Array_0_n1026, 
      load_n_store_RGB_Array_0_n1025, load_n_store_RGB_Array_0_n1024, 
      load_n_store_RGB_Array_0_n1023, load_n_store_RGB_Array_0_n1022, 
      load_n_store_RGB_Array_0_n1021, load_n_store_RGB_Array_0_n1020, 
      load_n_store_RGB_Array_0_n1019, load_n_store_RGB_Array_0_n1018, 
      load_n_store_RGB_Array_0_n1017, load_n_store_RGB_Array_0_n1016, 
      load_n_store_RGB_Array_0_n1015, load_n_store_RGB_Array_0_n1014, 
      load_n_store_RGB_Array_0_n1013, load_n_store_RGB_Array_0_n1012, 
      load_n_store_RGB_Array_0_n1011, load_n_store_RGB_Array_0_n1010, 
      load_n_store_RGB_Array_0_n1009, load_n_store_RGB_Array_0_n1008, 
      load_n_store_RGB_Array_0_n1007, load_n_store_RGB_Array_0_n1006, 
      load_n_store_RGB_Array_0_n1005, load_n_store_RGB_Array_0_n1004, 
      load_n_store_RGB_Array_0_n1003, load_n_store_RGB_Array_0_n1002, 
      load_n_store_RGB_Array_0_n1001, load_n_store_RGB_Array_0_n1000, 
      load_n_store_RGB_Array_0_n999, load_n_store_RGB_Array_0_n998, 
      load_n_store_RGB_Array_0_n997, load_n_store_RGB_Array_0_n996, 
      load_n_store_RGB_Array_0_n995, load_n_store_RGB_Array_0_n994, 
      load_n_store_RGB_Array_0_n993, load_n_store_RGB_Array_0_n992, 
      load_n_store_RGB_Array_0_n991, load_n_store_RGB_Array_0_n990, 
      load_n_store_RGB_Array_0_n989, load_n_store_RGB_Array_0_n988, 
      load_n_store_RGB_Array_0_n987, load_n_store_RGB_Array_0_n986, 
      load_n_store_RGB_Array_0_n985, load_n_store_RGB_Array_0_n984, 
      load_n_store_RGB_Array_0_n983, load_n_store_RGB_Array_0_n982, 
      load_n_store_RGB_Array_0_n981, load_n_store_RGB_Array_0_n980, 
      load_n_store_RGB_Array_0_n979, load_n_store_RGB_Array_0_n978, 
      load_n_store_RGB_Array_0_n977, load_n_store_RGB_Array_0_n976, 
      load_n_store_RGB_Array_0_n975, load_n_store_RGB_Array_0_n974, 
      load_n_store_RGB_Array_0_n973, load_n_store_RGB_Array_0_n972, 
      load_n_store_RGB_Array_0_n971, load_n_store_RGB_Array_0_n970, 
      load_n_store_RGB_Array_0_n969, load_n_store_RGB_Array_0_n968, 
      load_n_store_RGB_Array_0_n967, load_n_store_RGB_Array_0_n966, 
      load_n_store_RGB_Array_0_n965, load_n_store_RGB_Array_0_n964, 
      load_n_store_RGB_Array_0_n963, load_n_store_RGB_Array_0_n962, 
      load_n_store_RGB_Array_0_n961, load_n_store_RGB_Array_0_n960, 
      load_n_store_RGB_Array_0_n959, load_n_store_RGB_Array_0_n958, 
      load_n_store_RGB_Array_0_n957, load_n_store_RGB_Array_0_n956, 
      load_n_store_RGB_Array_0_n955, load_n_store_RGB_Array_0_n954, 
      load_n_store_RGB_Array_0_n953, load_n_store_RGB_Array_0_n952, 
      load_n_store_RGB_Array_0_n951, load_n_store_RGB_Array_0_n950, 
      load_n_store_RGB_Array_0_n949, load_n_store_RGB_Array_0_n948, 
      load_n_store_RGB_Array_0_n947, load_n_store_RGB_Array_0_n946, 
      load_n_store_RGB_Array_0_n945, load_n_store_RGB_Array_0_n944, 
      load_n_store_RGB_Array_0_n943, load_n_store_RGB_Array_0_n942, 
      load_n_store_RGB_Array_0_n941, load_n_store_RGB_Array_0_n940, 
      load_n_store_RGB_Array_0_n939, load_n_store_RGB_Array_0_n938, 
      load_n_store_RGB_Array_0_n937, load_n_store_RGB_Array_0_n936, 
      load_n_store_RGB_Array_0_n935, load_n_store_RGB_Array_0_n934, 
      load_n_store_RGB_Array_0_n933, load_n_store_RGB_Array_0_n932, 
      load_n_store_RGB_Array_0_n931, load_n_store_RGB_Array_0_n930, 
      load_n_store_RGB_Array_0_n929, load_n_store_RGB_Array_0_n928, 
      load_n_store_RGB_Array_0_n927, load_n_store_RGB_Array_0_n926, 
      load_n_store_RGB_Array_0_n925, load_n_store_RGB_Array_0_n924, 
      load_n_store_RGB_Array_0_n923, load_n_store_RGB_Array_0_n922, 
      load_n_store_RGB_Array_0_n921, load_n_store_RGB_Array_0_n920, 
      load_n_store_RGB_Array_0_n919, load_n_store_RGB_Array_0_n918, 
      load_n_store_RGB_Array_0_n917, load_n_store_RGB_Array_0_n916, 
      load_n_store_RGB_Array_0_n915, load_n_store_RGB_Array_0_n914, 
      load_n_store_RGB_Array_0_n913, load_n_store_RGB_Array_0_n912, 
      load_n_store_RGB_Array_0_n911, load_n_store_RGB_Array_0_n910, 
      load_n_store_RGB_Array_0_n909, load_n_store_RGB_Array_0_n908, 
      load_n_store_RGB_Array_0_n907, load_n_store_RGB_Array_0_n906, 
      load_n_store_RGB_Array_0_n905, load_n_store_RGB_Array_0_n904, 
      load_n_store_RGB_Array_0_n903, load_n_store_RGB_Array_0_n902, 
      load_n_store_RGB_Array_0_n901, load_n_store_RGB_Array_0_n900, 
      load_n_store_RGB_Array_0_n899, load_n_store_RGB_Array_0_n898, 
      load_n_store_RGB_Array_0_n897, load_n_store_RGB_Array_0_n896, 
      load_n_store_RGB_Array_0_n895, load_n_store_RGB_Array_0_n894, 
      load_n_store_RGB_Array_0_n893, load_n_store_RGB_Array_0_n892, 
      load_n_store_RGB_Array_0_n891, load_n_store_RGB_Array_0_n890, 
      load_n_store_RGB_Array_0_n889, load_n_store_RGB_Array_0_n888, 
      load_n_store_RGB_Array_0_n887, load_n_store_RGB_Array_0_n886, 
      load_n_store_RGB_Array_0_n885, load_n_store_RGB_Array_0_n884, 
      load_n_store_RGB_Array_0_n883, load_n_store_RGB_Array_0_n882, 
      load_n_store_RGB_Array_0_n881, load_n_store_RGB_Array_0_n880, 
      load_n_store_RGB_Array_0_n879, load_n_store_RGB_Array_0_n878, 
      load_n_store_RGB_Array_0_n877, load_n_store_RGB_Array_0_n876, 
      load_n_store_RGB_Array_0_n875, load_n_store_RGB_Array_0_n874, 
      load_n_store_RGB_Array_0_n873, load_n_store_RGB_Array_0_n872, 
      load_n_store_RGB_Array_0_n871, load_n_store_RGB_Array_0_n870, 
      load_n_store_RGB_Array_0_n869, load_n_store_RGB_Array_0_n868, 
      load_n_store_RGB_Array_0_n867, load_n_store_RGB_Array_0_n866, 
      load_n_store_RGB_Array_0_n865, load_n_store_RGB_Array_0_n864, 
      load_n_store_RGB_Array_0_n863, load_n_store_RGB_Array_0_n862, 
      load_n_store_RGB_Array_0_n861, load_n_store_RGB_Array_0_n860, 
      load_n_store_RGB_Array_0_n859, load_n_store_RGB_Array_0_n858, 
      load_n_store_RGB_Array_0_n857, load_n_store_RGB_Array_0_n856, 
      load_n_store_RGB_Array_0_n855, load_n_store_RGB_Array_0_n854, 
      load_n_store_RGB_Array_0_n853, load_n_store_RGB_Array_0_n852, 
      load_n_store_RGB_Array_0_n851, load_n_store_RGB_Array_0_n850, 
      load_n_store_RGB_Array_0_n849, load_n_store_RGB_Array_0_n848, 
      load_n_store_RGB_Array_0_n847, load_n_store_RGB_Array_0_n846, 
      load_n_store_RGB_Array_0_n845, load_n_store_RGB_Array_0_n844, 
      load_n_store_RGB_Array_0_n843, load_n_store_RGB_Array_0_n842, 
      load_n_store_RGB_Array_0_n841, load_n_store_RGB_Array_0_n840, 
      load_n_store_RGB_Array_0_n839, load_n_store_RGB_Array_0_n838, 
      load_n_store_RGB_Array_0_n837, load_n_store_RGB_Array_0_n836, 
      load_n_store_RGB_Array_0_n835, load_n_store_RGB_Array_0_n834, 
      load_n_store_RGB_Array_0_n833, load_n_store_RGB_Array_0_n832, 
      load_n_store_RGB_Array_0_n831, load_n_store_RGB_Array_0_n830, 
      load_n_store_RGB_Array_0_n829, load_n_store_RGB_Array_0_n828, 
      load_n_store_RGB_Array_0_n827, load_n_store_RGB_Array_0_n826, 
      load_n_store_RGB_Array_0_n825, load_n_store_RGB_Array_0_n824, 
      load_n_store_RGB_Array_0_n823, load_n_store_RGB_Array_0_n822, 
      load_n_store_RGB_Array_0_n821, load_n_store_RGB_Array_0_n820, 
      load_n_store_RGB_Array_0_n819, load_n_store_RGB_Array_0_n818, 
      load_n_store_RGB_Array_0_n817, load_n_store_RGB_Array_0_n816, 
      load_n_store_RGB_Array_0_n815, load_n_store_RGB_Array_0_n814, 
      load_n_store_RGB_Array_0_n813, load_n_store_RGB_Array_0_n812, 
      load_n_store_RGB_Array_0_n811, load_n_store_RGB_Array_0_n810, 
      load_n_store_RGB_Array_0_n809, load_n_store_RGB_Array_0_n808, 
      load_n_store_RGB_Array_0_n807, load_n_store_RGB_Array_0_n806, 
      load_n_store_RGB_Array_0_n805, load_n_store_RGB_Array_0_n804, 
      load_n_store_RGB_Array_0_n803, load_n_store_RGB_Array_0_n802, 
      load_n_store_RGB_Array_0_n801, load_n_store_RGB_Array_0_n800, 
      load_n_store_RGB_Array_0_n799, load_n_store_RGB_Array_0_n798, 
      load_n_store_RGB_Array_0_n797, load_n_store_RGB_Array_0_n796, 
      load_n_store_RGB_Array_0_n795, load_n_store_RGB_Array_0_n794, 
      load_n_store_RGB_Array_0_n793, load_n_store_RGB_Array_0_n792, 
      load_n_store_RGB_Array_0_n791, load_n_store_RGB_Array_0_n790, 
      load_n_store_RGB_Array_0_n789, load_n_store_RGB_Array_0_n788, 
      load_n_store_RGB_Array_0_n787, load_n_store_RGB_Array_0_n786, 
      load_n_store_RGB_Array_0_n785, load_n_store_RGB_Array_0_n784, 
      load_n_store_RGB_Array_0_n783, load_n_store_RGB_Array_0_n782, 
      load_n_store_RGB_Array_0_n781, load_n_store_RGB_Array_0_n780, 
      load_n_store_RGB_Array_0_n779, load_n_store_RGB_Array_0_n778, 
      load_n_store_RGB_Array_0_n777, load_n_store_RGB_Array_0_n776, 
      load_n_store_RGB_Array_0_n775, load_n_store_RGB_Array_0_n774, 
      load_n_store_RGB_Array_0_n773, load_n_store_RGB_Array_0_n772, 
      load_n_store_RGB_Array_0_n771, load_n_store_RGB_Array_0_n770, 
      load_n_store_RGB_Array_0_n769, load_n_store_RGB_Array_0_n768, 
      load_n_store_RGB_Array_0_n767, load_n_store_RGB_Array_0_n766, 
      load_n_store_RGB_Array_0_n765, load_n_store_RGB_Array_0_n764, 
      load_n_store_RGB_Array_0_n763, load_n_store_RGB_Array_0_n762, 
      load_n_store_RGB_Array_0_n761, load_n_store_RGB_Array_0_n760, 
      load_n_store_RGB_Array_0_n759, load_n_store_RGB_Array_0_n758, 
      load_n_store_RGB_Array_0_n757, load_n_store_RGB_Array_0_n756, 
      load_n_store_RGB_Array_0_n755, load_n_store_RGB_Array_0_n754, 
      load_n_store_RGB_Array_0_n753, load_n_store_RGB_Array_0_n752, 
      load_n_store_RGB_Array_0_n751, load_n_store_RGB_Array_0_n750, 
      load_n_store_RGB_Array_0_n749, load_n_store_RGB_Array_0_n748, 
      load_n_store_RGB_Array_0_n747, load_n_store_RGB_Array_0_n746, 
      load_n_store_RGB_Array_0_n745, load_n_store_RGB_Array_0_n744, 
      load_n_store_RGB_Array_0_n743, load_n_store_RGB_Array_0_n742, 
      load_n_store_RGB_Array_0_n741, load_n_store_RGB_Array_0_n740, 
      load_n_store_RGB_Array_0_n739, load_n_store_RGB_Array_0_n738, 
      load_n_store_RGB_Array_0_n737, load_n_store_RGB_Array_0_n736, 
      load_n_store_RGB_Array_0_n735, load_n_store_RGB_Array_0_n734, 
      load_n_store_RGB_Array_0_n733, load_n_store_RGB_Array_0_n732, 
      load_n_store_RGB_Array_0_n731, load_n_store_RGB_Array_0_n730, 
      load_n_store_RGB_Array_0_n729, load_n_store_RGB_Array_0_n728, 
      load_n_store_RGB_Array_0_n727, load_n_store_RGB_Array_0_n726, 
      load_n_store_RGB_Array_0_n725, load_n_store_RGB_Array_0_n724, 
      load_n_store_RGB_Array_0_n723, load_n_store_RGB_Array_0_n722, 
      load_n_store_RGB_Array_0_n721, load_n_store_RGB_Array_0_n720, 
      load_n_store_RGB_Array_0_n719, load_n_store_RGB_Array_0_n718, 
      load_n_store_RGB_Array_0_n717, load_n_store_RGB_Array_0_n716, 
      load_n_store_RGB_Array_0_n715, load_n_store_RGB_Array_0_n714, 
      load_n_store_RGB_Array_0_n713, load_n_store_RGB_Array_0_n712, 
      load_n_store_RGB_Array_0_n711, load_n_store_RGB_Array_0_n710, 
      load_n_store_RGB_Array_0_n709, load_n_store_RGB_Array_0_n708, 
      load_n_store_RGB_Array_0_n707, load_n_store_RGB_Array_0_n706, 
      load_n_store_RGB_Array_0_n705, load_n_store_RGB_Array_0_n704, 
      load_n_store_RGB_Array_0_n703, load_n_store_RGB_Array_0_n702, 
      load_n_store_RGB_Array_0_n701, load_n_store_RGB_Array_0_n700, 
      load_n_store_RGB_Array_0_n699, load_n_store_RGB_Array_0_n698, 
      load_n_store_RGB_Array_0_n697, load_n_store_RGB_Array_0_n696, 
      load_n_store_RGB_Array_0_n695, load_n_store_RGB_Array_0_n694, 
      load_n_store_RGB_Array_0_n693, load_n_store_RGB_Array_0_n692, 
      load_n_store_RGB_Array_0_n691, load_n_store_RGB_Array_0_n690, 
      load_n_store_RGB_Array_0_n689, load_n_store_RGB_Array_0_n688, 
      load_n_store_RGB_Array_0_n687, load_n_store_RGB_Array_0_n686, 
      load_n_store_RGB_Array_0_n685, load_n_store_RGB_Array_0_n684, 
      load_n_store_RGB_Array_0_n683, load_n_store_RGB_Array_0_n682, 
      load_n_store_RGB_Array_0_n681, load_n_store_RGB_Array_0_n680, 
      load_n_store_RGB_Array_0_n679, load_n_store_RGB_Array_0_n678, 
      load_n_store_RGB_Array_0_n677, load_n_store_RGB_Array_0_n676, 
      load_n_store_RGB_Array_0_n675, load_n_store_RGB_Array_0_n674, 
      load_n_store_RGB_Array_0_n673, load_n_store_RGB_Array_0_n672, 
      load_n_store_RGB_Array_0_n671, load_n_store_RGB_Array_0_n670, 
      load_n_store_RGB_Array_0_n669, load_n_store_RGB_Array_0_n668, 
      load_n_store_RGB_Array_0_n667, load_n_store_RGB_Array_0_n666, 
      load_n_store_RGB_Array_0_n665, load_n_store_RGB_Array_0_n664, 
      load_n_store_RGB_Array_0_n663, load_n_store_RGB_Array_0_n662, 
      load_n_store_RGB_Array_0_n661, load_n_store_RGB_Array_0_n660, 
      load_n_store_RGB_Array_0_n659, load_n_store_RGB_Array_0_n658, 
      load_n_store_RGB_Array_0_n657, load_n_store_RGB_Array_0_n656, 
      load_n_store_RGB_Array_0_n655, load_n_store_RGB_Array_0_n654, 
      load_n_store_RGB_Array_0_n653, load_n_store_RGB_Array_0_n652, 
      load_n_store_RGB_Array_0_n651, load_n_store_RGB_Array_0_n650, 
      load_n_store_RGB_Array_0_n649, load_n_store_RGB_Array_0_n648, 
      load_n_store_RGB_Array_0_n647, load_n_store_RGB_Array_0_n646, 
      load_n_store_RGB_Array_0_n645, load_n_store_RGB_Array_0_n644, 
      load_n_store_RGB_Array_0_n643, load_n_store_RGB_Array_0_n642, 
      load_n_store_RGB_Array_0_n641, load_n_store_RGB_Array_0_n640, 
      load_n_store_RGB_Array_0_n639, load_n_store_RGB_Array_0_n638, 
      load_n_store_RGB_Array_0_n637, load_n_store_RGB_Array_0_n636, 
      load_n_store_RGB_Array_0_n635, 
      load_n_store_RGB_Array_0_block_ram_r_0_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_0_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_0_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_0_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_0_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_0_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_0_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_0_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_1_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_1_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_1_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_1_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_1_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_1_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_1_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_1_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_2_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_2_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_2_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_2_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_2_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_2_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_2_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_2_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_3_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_3_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_3_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_3_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_3_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_3_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_3_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_3_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_4_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_4_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_4_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_4_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_4_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_4_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_4_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_4_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_5_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_5_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_5_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_5_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_5_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_5_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_5_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_5_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_6_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_6_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_6_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_6_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_6_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_6_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_6_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_6_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_7_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_7_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_7_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_7_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_7_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_7_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_7_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_7_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_8_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_8_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_8_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_8_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_8_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_8_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_8_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_8_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_9_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_9_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_9_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_9_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_9_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_9_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_9_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_9_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_10_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_10_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_10_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_10_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_10_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_10_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_10_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_10_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_11_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_11_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_11_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_11_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_11_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_11_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_11_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_11_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_12_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_12_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_12_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_12_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_12_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_12_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_12_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_12_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_13_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_13_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_13_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_13_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_13_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_13_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_13_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_13_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_14_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_14_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_14_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_14_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_14_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_14_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_14_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_14_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_15_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_15_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_15_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_15_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_15_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_15_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_15_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_15_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_16_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_16_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_16_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_16_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_16_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_16_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_16_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_16_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_17_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_17_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_17_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_17_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_17_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_17_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_17_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_17_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_18_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_18_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_18_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_18_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_18_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_18_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_18_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_18_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_19_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_19_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_19_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_19_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_19_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_19_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_19_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_19_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_20_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_20_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_20_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_20_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_20_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_20_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_20_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_20_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_21_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_21_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_21_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_21_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_21_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_21_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_21_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_21_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_22_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_22_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_22_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_22_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_22_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_22_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_22_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_22_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_23_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_23_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_23_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_23_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_23_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_23_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_23_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_23_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_24_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_24_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_24_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_24_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_24_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_24_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_24_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_24_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_25_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_25_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_25_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_25_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_25_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_25_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_25_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_25_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_26_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_26_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_26_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_26_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_26_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_26_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_26_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_26_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_27_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_27_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_27_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_27_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_27_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_27_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_27_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_27_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_28_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_28_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_28_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_28_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_28_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_28_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_28_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_28_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_29_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_29_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_29_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_29_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_29_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_29_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_29_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_29_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_30_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_30_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_30_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_30_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_30_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_30_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_30_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_30_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_31_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_31_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_31_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_31_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_31_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_31_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_31_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_31_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_0_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_0_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_0_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_0_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_0_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_0_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_0_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_0_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_1_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_1_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_1_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_1_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_1_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_1_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_1_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_1_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_2_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_2_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_2_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_2_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_2_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_2_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_2_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_2_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_3_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_3_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_3_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_3_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_3_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_3_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_3_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_3_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_4_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_4_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_4_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_4_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_4_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_4_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_4_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_4_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_5_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_5_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_5_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_5_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_5_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_5_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_5_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_5_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_6_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_6_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_6_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_6_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_6_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_6_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_6_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_6_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_7_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_7_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_7_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_7_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_7_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_7_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_7_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_7_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_8_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_8_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_8_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_8_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_8_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_8_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_8_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_8_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_9_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_9_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_9_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_9_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_9_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_9_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_9_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_9_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_10_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_10_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_10_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_10_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_10_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_10_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_10_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_10_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_11_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_11_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_11_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_11_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_11_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_11_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_11_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_11_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_12_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_12_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_12_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_12_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_12_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_12_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_12_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_12_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_13_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_13_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_13_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_13_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_13_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_13_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_13_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_13_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_14_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_14_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_14_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_14_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_14_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_14_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_14_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_14_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_15_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_15_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_15_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_15_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_15_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_15_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_15_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_15_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_16_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_16_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_16_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_16_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_16_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_16_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_16_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_16_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_17_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_17_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_17_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_17_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_17_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_17_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_17_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_17_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_18_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_18_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_18_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_18_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_18_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_18_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_18_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_18_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_19_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_19_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_19_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_19_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_19_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_19_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_19_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_19_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_20_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_20_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_20_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_20_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_20_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_20_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_20_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_20_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_21_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_21_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_21_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_21_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_21_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_21_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_21_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_21_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_22_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_22_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_22_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_22_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_22_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_22_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_22_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_22_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_23_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_23_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_23_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_23_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_23_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_23_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_23_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_23_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_24_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_24_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_24_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_24_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_24_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_24_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_24_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_24_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_25_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_25_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_25_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_25_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_25_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_25_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_25_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_25_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_26_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_26_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_26_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_26_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_26_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_26_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_26_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_26_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_27_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_27_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_27_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_27_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_27_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_27_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_27_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_27_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_28_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_28_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_28_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_28_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_28_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_28_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_28_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_28_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_29_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_29_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_29_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_29_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_29_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_29_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_29_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_29_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_30_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_30_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_30_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_30_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_30_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_30_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_30_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_30_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_31_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_31_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_31_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_31_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_31_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_31_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_31_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_31_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_0_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_0_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_0_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_0_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_0_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_0_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_0_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_0_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_1_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_1_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_1_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_1_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_1_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_1_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_1_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_1_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_2_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_2_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_2_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_2_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_2_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_2_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_2_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_2_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_3_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_3_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_3_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_3_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_3_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_3_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_3_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_3_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_4_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_4_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_4_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_4_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_4_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_4_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_4_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_4_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_5_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_5_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_5_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_5_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_5_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_5_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_5_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_5_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_6_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_6_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_6_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_6_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_6_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_6_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_6_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_6_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_7_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_7_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_7_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_7_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_7_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_7_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_7_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_7_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_8_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_8_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_8_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_8_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_8_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_8_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_8_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_8_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_9_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_9_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_9_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_9_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_9_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_9_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_9_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_9_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_10_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_10_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_10_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_10_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_10_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_10_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_10_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_10_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_11_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_11_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_11_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_11_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_11_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_11_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_11_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_11_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_12_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_12_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_12_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_12_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_12_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_12_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_12_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_12_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_13_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_13_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_13_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_13_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_13_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_13_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_13_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_13_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_14_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_14_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_14_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_14_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_14_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_14_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_14_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_14_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_15_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_15_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_15_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_15_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_15_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_15_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_15_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_15_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_16_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_16_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_16_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_16_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_16_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_16_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_16_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_16_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_17_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_17_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_17_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_17_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_17_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_17_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_17_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_17_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_18_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_18_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_18_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_18_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_18_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_18_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_18_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_18_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_19_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_19_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_19_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_19_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_19_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_19_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_19_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_19_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_20_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_20_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_20_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_20_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_20_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_20_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_20_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_20_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_21_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_21_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_21_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_21_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_21_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_21_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_21_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_21_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_22_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_22_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_22_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_22_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_22_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_22_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_22_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_22_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_23_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_23_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_23_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_23_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_23_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_23_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_23_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_23_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_24_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_24_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_24_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_24_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_24_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_24_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_24_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_24_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_25_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_25_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_25_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_25_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_25_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_25_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_25_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_25_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_26_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_26_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_26_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_26_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_26_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_26_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_26_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_26_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_27_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_27_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_27_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_27_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_27_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_27_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_27_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_27_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_28_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_28_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_28_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_28_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_28_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_28_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_28_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_28_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_29_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_29_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_29_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_29_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_29_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_29_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_29_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_29_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_30_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_30_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_30_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_30_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_30_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_30_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_30_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_30_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_31_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_31_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_31_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_31_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_31_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_31_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_31_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_31_7_port, n1, n2, n3, n4, n5, n6, 
      n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
      n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
      n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, 
      n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
      n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, 
      n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, 
      n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, 
      n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, 
      n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, 
      n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, 
      n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, 
      n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, 
      n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, 
      n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, 
      n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, 
      n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, 
      n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, 
      n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, 
      n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, 
      n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, 
      n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, 
      n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, 
      n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, 
      n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, 
      n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, 
      n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, 
      n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, 
      n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, 
      n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, 
      n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, 
      n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, 
      n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, 
      n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, 
      n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, 
      n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, 
      n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, 
      n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, 
      n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, 
      n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, 
      n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, 
      n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, 
      n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, 
      n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, 
      n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, 
      n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, 
      n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, 
      n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, 
      n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, 
      n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, 
      n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, 
      n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, 
      n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, 
      n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, 
      n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, 
      n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, 
      n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, 
      n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, 
      n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, 
      n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, 
      n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, 
      n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, 
      n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, 
      n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, 
      n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, 
      n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, 
      n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, 
      n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, 
      n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, 
      n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, 
      n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, 
      n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, 
      n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, 
      n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, 
      n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, 
      n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, 
      n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, 
      n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, 
      n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, 
      n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, 
      n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
      n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, 
      n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, 
      n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, 
      n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, 
      n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, 
      n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
      n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
      n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
      n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
      n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, 
      n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
      n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, 
      n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, 
      n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
      n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
      n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
      n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
      n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
      n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
      n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
      n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
      n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, 
      n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
      n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
      n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, 
      n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, 
      n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, 
      n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, 
      n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, 
      n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, 
      n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, 
      n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, 
      n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, 
      n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, 
      n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, 
      n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, 
      n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, 
      n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, 
      n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, 
      n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, 
      n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, 
      n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, 
      n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, 
      n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, 
      n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, 
      n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, 
      n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
      n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, 
      n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, 
      n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, 
      n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, 
      n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, 
      n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, 
      n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, 
      n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, 
      n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, 
      n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, 
      n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, 
      n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, 
      n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, 
      n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, 
      n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, 
      n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, 
      n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, 
      n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, 
      n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, 
      n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, 
      n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, 
      n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, 
      n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, 
      n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, 
      n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, 
      n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, 
      n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, 
      n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, 
      n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, 
      n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, 
      n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, 
      n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, 
      n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, 
      n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, 
      n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, 
      n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, 
      n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, 
      n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, 
      n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, 
      n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, 
      n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, 
      n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, 
      n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, 
      n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, 
      n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, 
      n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, 
      n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, 
      n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, 
      n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, 
      n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, 
      n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, 
      n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, 
      n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, 
      n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, 
      n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, 
      n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, 
      n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, 
      n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, 
      n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, 
      n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, 
      n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, 
      n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, 
      n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, 
      n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, 
      n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, 
      n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, 
      n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, 
      n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, 
      n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, 
      n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, 
      n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, 
      n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, 
      n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, 
      n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, 
      n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, 
      n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, 
      n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, 
      n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, 
      n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, 
      n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, 
      n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, 
      n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, 
      n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, 
      n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, 
      n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, 
      n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, 
      n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, 
      n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, 
      n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, 
      n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, 
      n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, 
      n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, 
      n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, 
      n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, 
      n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344 : bit;

begin
   reset_port <= reset;
   top_ack <= top_ack_port;
   hub_mux_o <= ( hub_mux_o_2_port, hub_mux_o_1_port, hub_mux_o_0_port );
   hub_clk_o <= hub_clk_o_port;
   hub_latch_o <= hub_latch_o_port;
   hub_blank_o <= hub_blank_o_port;
   hub_g0_o <= hub_g0_o_port;
   hub_b0_o <= hub_b0_o_port;
   hub_r0_o <= hub_r0_o_port;
   
   registers_n84 <= '1';
   registers_n83 <= '1';
   registers_n82 <= '1';
   registers_n81 <= '1';
   registers_n80 <= '1';
   registers_n79 <= '1';
   registers_n78 <= '1';
   registers_n77 <= '1';
   registers_n76 <= '1';
   registers_n75 <= '1';
   registers_n74 <= '1';
   registers_n73 <= '1';
   registers_n72 <= '1';
   registers_n71 <= '1';
   registers_n70 <= '1';
   registers_n69 <= '1';
   registers_n68 <= '1';
   registers_n67 <= '1';
   registers_n66 <= '1';
   registers_n65 <= '1';
   registers_n64 <= '1';
   registers_n63 <= '1';
   registers_n62 <= '1';
   registers_n61 <= '1';
   registers_n60 <= '1';
   registers_n59 <= '1';
   registers_n58 <= '1';
   registers_n57 <= '1';
   registers_n56 <= '1';
   registers_n55 <= '1';
   registers_n54 <= '1';
   registers_n53 <= '1';
   registers_n52 <= '1';
   registers_n51 <= '1';
   registers_n50 <= '1';
   registers_n49 <= '1';
   registers_n48 <= '1';
   registers_n47 <= '1';
   registers_n46 <= '1';
   registers_n45 <= '1';
   registers_n44 <= '1';
   registers_n43 <= '1';
   registers_n42 <= '1';
   registers_n41 <= '1';
   registers_n40 <= '1';
   registers_n39 <= '1';
   registers_n38 <= '1';
   registers_n37 <= '1';
   registers_n36 <= '1';
   registers_n35 <= '1';
   registers_n34 <= '1';
   registers_n33 <= '1';
   registers_n32 <= '1';
   registers_n31 <= '1';
   registers_n30 <= '1';
   registers_n29 <= '1';
   registers_n28 <= '1';
   registers_n27 <= '1';
   registers_n26 <= '1';
   registers_n25 <= '1';
   registers_n24 <= '1';
   registers_n23 <= '1';
   registers_n22 <= '1';
   registers_n21 <= '1';
   registers_n20 <= '1';
   registers_n19 <= '1';
   registers_mem_sipo_g0_reg_0_inst : dff port map( d => registers_n232, gclk 
                           => clk, rnot => registers_n19, q => 
                           mem_sipo_g0_0_port);
   registers_mem_sipo_g0_reg_1_inst : dff port map( d => registers_n233, gclk 
                           => clk, rnot => registers_n20, q => 
                           mem_sipo_g0_1_port);
   registers_mem_sipo_g0_reg_2_inst : dff port map( d => registers_n234, gclk 
                           => clk, rnot => registers_n21, q => 
                           mem_sipo_g0_2_port);
   registers_mem_sipo_g0_reg_3_inst : dff port map( d => registers_n235, gclk 
                           => clk, rnot => registers_n22, q => 
                           mem_sipo_g0_3_port);
   registers_mem_sipo_g0_reg_4_inst : dff port map( d => registers_n236, gclk 
                           => clk, rnot => registers_n23, q => 
                           mem_sipo_g0_4_port);
   registers_mem_sipo_g0_reg_5_inst : dff port map( d => registers_n237, gclk 
                           => clk, rnot => registers_n24, q => 
                           mem_sipo_g0_5_port);
   registers_mem_sipo_g0_reg_6_inst : dff port map( d => registers_n238, gclk 
                           => clk, rnot => registers_n25, q => 
                           mem_sipo_g0_6_port);
   registers_mem_sipo_g0_reg_7_inst : dff port map( d => registers_n239, gclk 
                           => clk, rnot => registers_n26, q => 
                           mem_sipo_g0_7_port);
   registers_mem_sipo_r0_reg_0_inst : dff port map( d => registers_n240, gclk 
                           => clk, rnot => registers_n27, q => 
                           mem_sipo_r0_0_port);
   registers_mem_sipo_r0_reg_1_inst : dff port map( d => registers_n241, gclk 
                           => clk, rnot => registers_n28, q => 
                           mem_sipo_r0_1_port);
   registers_mem_sipo_r0_reg_2_inst : dff port map( d => registers_n242, gclk 
                           => clk, rnot => registers_n29, q => 
                           mem_sipo_r0_2_port);
   registers_mem_sipo_r0_reg_3_inst : dff port map( d => registers_n243, gclk 
                           => clk, rnot => registers_n30, q => 
                           mem_sipo_r0_3_port);
   registers_mem_sipo_r0_reg_4_inst : dff port map( d => registers_n244, gclk 
                           => clk, rnot => registers_n31, q => 
                           mem_sipo_r0_4_port);
   registers_mem_sipo_r0_reg_5_inst : dff port map( d => registers_n245, gclk 
                           => clk, rnot => registers_n32, q => 
                           mem_sipo_r0_5_port);
   registers_mem_sipo_r0_reg_6_inst : dff port map( d => registers_n246, gclk 
                           => clk, rnot => registers_n33, q => 
                           mem_sipo_r0_6_port);
   registers_mem_sipo_r0_reg_7_inst : dff port map( d => registers_n247, gclk 
                           => clk, rnot => registers_n34, q => 
                           mem_sipo_r0_7_port);
   registers_s_mem_sipo_g0_reg_0_inst : dff port map( d => registers_n248, gclk
                           => clk, rnot => registers_n35, q => 
                           registers_s_mem_sipo_g0_0_port);
   registers_s_mem_sipo_g0_reg_1_inst : dff port map( d => registers_n249, gclk
                           => clk, rnot => registers_n36, q => 
                           registers_s_mem_sipo_g0_1_port);
   registers_s_mem_sipo_g0_reg_2_inst : dff port map( d => registers_n250, gclk
                           => clk, rnot => registers_n37, q => 
                           registers_s_mem_sipo_g0_2_port);
   registers_s_mem_sipo_g0_reg_3_inst : dff port map( d => registers_n251, gclk
                           => clk, rnot => registers_n38, q => 
                           registers_s_mem_sipo_g0_3_port);
   registers_s_mem_sipo_g0_reg_4_inst : dff port map( d => registers_n252, gclk
                           => clk, rnot => registers_n39, q => 
                           registers_s_mem_sipo_g0_4_port);
   registers_s_mem_sipo_g0_reg_5_inst : dff port map( d => registers_n253, gclk
                           => clk, rnot => registers_n40, q => 
                           registers_s_mem_sipo_g0_5_port);
   registers_s_mem_sipo_g0_reg_6_inst : dff port map( d => registers_n254, gclk
                           => clk, rnot => registers_n41, q => 
                           registers_s_mem_sipo_g0_6_port);
   registers_s_mem_sipo_g0_reg_7_inst : dff port map( d => registers_n255, gclk
                           => clk, rnot => registers_n42, q => 
                           registers_s_mem_sipo_g0_7_port);
   registers_s_mem_sipo_r0_reg_0_inst : dff port map( d => registers_n256, gclk
                           => clk, rnot => registers_n43, q => 
                           registers_s_mem_sipo_r0_0_port);
   registers_s_mem_sipo_r0_reg_1_inst : dff port map( d => registers_n257, gclk
                           => clk, rnot => registers_n44, q => 
                           registers_s_mem_sipo_r0_1_port);
   registers_s_mem_sipo_r0_reg_2_inst : dff port map( d => registers_n258, gclk
                           => clk, rnot => registers_n45, q => 
                           registers_s_mem_sipo_r0_2_port);
   registers_s_mem_sipo_r0_reg_3_inst : dff port map( d => registers_n259, gclk
                           => clk, rnot => registers_n46, q => 
                           registers_s_mem_sipo_r0_3_port);
   registers_s_mem_sipo_r0_reg_4_inst : dff port map( d => registers_n260, gclk
                           => clk, rnot => registers_n47, q => 
                           registers_s_mem_sipo_r0_4_port);
   registers_s_mem_sipo_r0_reg_5_inst : dff port map( d => registers_n261, gclk
                           => clk, rnot => registers_n48, q => 
                           registers_s_mem_sipo_r0_5_port);
   registers_s_mem_sipo_r0_reg_6_inst : dff port map( d => registers_n262, gclk
                           => clk, rnot => registers_n49, q => 
                           registers_s_mem_sipo_r0_6_port);
   registers_s_mem_sipo_r0_reg_7_inst : dff port map( d => registers_n263, gclk
                           => clk, rnot => registers_n50, q => 
                           registers_s_mem_sipo_r0_7_port);
   registers_mem_sipo_b0_reg_0_inst : dff port map( d => registers_n264, gclk 
                           => clk, rnot => registers_n51, q => 
                           mem_sipo_b0_0_port);
   registers_s_mem_sipo_b0_reg_0_inst : dff port map( d => registers_n265, gclk
                           => clk, rnot => registers_n52, q => 
                           registers_s_mem_sipo_b0_0_port);
   registers_mem_sipo_b0_reg_1_inst : dff port map( d => registers_n266, gclk 
                           => clk, rnot => registers_n53, q => 
                           mem_sipo_b0_1_port);
   registers_s_mem_sipo_b0_reg_1_inst : dff port map( d => registers_n267, gclk
                           => clk, rnot => registers_n54, q => 
                           registers_s_mem_sipo_b0_1_port);
   registers_mem_sipo_b0_reg_2_inst : dff port map( d => registers_n268, gclk 
                           => clk, rnot => registers_n55, q => 
                           mem_sipo_b0_2_port);
   registers_s_mem_sipo_b0_reg_2_inst : dff port map( d => registers_n269, gclk
                           => clk, rnot => registers_n56, q => 
                           registers_s_mem_sipo_b0_2_port);
   registers_mem_sipo_b0_reg_3_inst : dff port map( d => registers_n270, gclk 
                           => clk, rnot => registers_n57, q => 
                           mem_sipo_b0_3_port);
   registers_s_mem_sipo_b0_reg_3_inst : dff port map( d => registers_n271, gclk
                           => clk, rnot => registers_n58, q => 
                           registers_s_mem_sipo_b0_3_port);
   registers_mem_sipo_b0_reg_4_inst : dff port map( d => registers_n272, gclk 
                           => clk, rnot => registers_n59, q => 
                           mem_sipo_b0_4_port);
   registers_s_mem_sipo_b0_reg_4_inst : dff port map( d => registers_n273, gclk
                           => clk, rnot => registers_n60, q => 
                           registers_s_mem_sipo_b0_4_port);
   registers_mem_sipo_b0_reg_5_inst : dff port map( d => registers_n274, gclk 
                           => clk, rnot => registers_n61, q => 
                           mem_sipo_b0_5_port);
   registers_s_mem_sipo_b0_reg_5_inst : dff port map( d => registers_n275, gclk
                           => clk, rnot => registers_n62, q => 
                           registers_s_mem_sipo_b0_5_port);
   registers_mem_sipo_b0_reg_6_inst : dff port map( d => registers_n276, gclk 
                           => clk, rnot => registers_n63, q => 
                           mem_sipo_b0_6_port);
   registers_s_mem_sipo_b0_reg_6_inst : dff port map( d => registers_n277, gclk
                           => clk, rnot => registers_n64, q => 
                           registers_s_mem_sipo_b0_6_port);
   registers_mem_sipo_b0_reg_7_inst : dff port map( d => registers_n278, gclk 
                           => clk, rnot => registers_n65, q => 
                           mem_sipo_b0_7_port);
   registers_s_mem_sipo_b0_reg_7_inst : dff port map( d => registers_n279, gclk
                           => clk, rnot => registers_n66, q => 
                           registers_s_mem_sipo_b0_7_port);
   registers_reg_hub_f_reg : dff port map( d => registers_n280, gclk => clk, 
                           rnot => registers_n67, q => reg_hub_f);
   registers_addr_i_reg_1_inst : dff port map( d => registers_n288, gclk => clk
                           , rnot => registers_n68, q => addr_i_1_port);
   registers_addr_i_reg_2_inst : dff port map( d => registers_n292, gclk => clk
                           , rnot => registers_n69, q => addr_i_2_port);
   registers_addr_i_reg_0_inst : dff port map( d => registers_n290, gclk => clk
                           , rnot => registers_n70, q => addr_i_0_port);
   registers_addr_i_reg_4_inst : dff port map( d => registers_n283, gclk => clk
                           , rnot => registers_n71, q => addr_i_4_port);
   registers_addr_i_reg_3_inst : dff port map( d => registers_n281, gclk => clk
                           , rnot => registers_n72, q => addr_i_3_port);
   registers_reg_row_reg_1_inst : dff port map( d => registers_n284, gclk => 
                           clk, rnot => registers_n73, q => 
                           registers_reg_row_1_port);
   registers_reg_cd_reg_0_inst : dff port map( d => registers_n286, gclk => clk
                           , rnot => registers_n74, q => 
                           registers_reg_cd_0_port);
   registers_reg_cd_reg_2_inst : dff port map( d => registers_n287, gclk => clk
                           , rnot => registers_n75, q => 
                           registers_reg_cd_2_port);
   registers_reg_cd_reg_1_inst : dff port map( d => registers_n285, gclk => clk
                           , rnot => registers_n76, q => 
                           registers_reg_cd_1_port);
   registers_reg_row_reg_0_inst : dff port map( d => registers_n282, gclk => 
                           clk, rnot => registers_n77, q => 
                           registers_reg_row_0_port);
   registers_mem_to_reg_reg_1_inst : dff port map( d => registers_n294, gclk =>
                           clk, rnot => registers_n78, q => 
                           registers_mem_to_reg_1_port);
   registers_reg_col_inc_reg_2_inst : dff port map( d => registers_n293, gclk 
                           => clk, rnot => registers_n79, q => 
                           registers_reg_col_inc_2_port);
   registers_reg_col_inc_reg_0_inst : dff port map( d => registers_n291, gclk 
                           => clk, rnot => registers_n80, q => 
                           registers_reg_col_inc_0_port);
   registers_reg_col_inc_reg_1_inst : dff port map( d => registers_n289, gclk 
                           => clk, rnot => registers_n81, q => 
                           registers_reg_col_inc_1_port);
   registers_mem_to_reg_reg_0_inst : dff port map( d => n2272, gclk => clk, 
                           rnot => registers_n82, q => 
                           registers_mem_to_reg_0_port);
   registers_s_delay_reg_1_inst : dff port map( d => registers_n295, gclk => 
                           clk, rnot => registers_n83, q => 
                           registers_s_delay_1_port);
   registers_s_delay_reg_0_inst : dff port map( d => registers_n296, gclk => 
                           clk, rnot => registers_n84, q => 
                           registers_s_delay_0_port);
   load_n_store_n76 <= '1';
   load_n_store_n75 <= '1';
   load_n_store_n74 <= '1';
   load_n_store_n73 <= '1';
   load_n_store_n72 <= '1';
   load_n_store_n71 <= '1';
   load_n_store_n70 <= '1';
   load_n_store_n69 <= '1';
   load_n_store_n68 <= '1';
   load_n_store_n67 <= '1';
   load_n_store_n66 <= '1';
   load_n_store_n65 <= '1';
   load_n_store_n64 <= '1';
   load_n_store_n63 <= '1';
   load_n_store_n62 <= '1';
   load_n_store_n61 <= '1';
   load_n_store_n60 <= '1';
   load_n_store_n59 <= '1';
   load_n_store_n58 <= '1';
   load_n_store_n57 <= '1';
   load_n_store_n56 <= '1';
   load_n_store_n55 <= '1';
   load_n_store_n54 <= '1';
   load_n_store_n53 <= '1';
   load_n_store_n52 <= '1';
   load_n_store_n51 <= '1';
   load_n_store_n50 <= '1';
   load_n_store_n49 <= '1';
   load_n_store_n48 <= '1';
   load_n_store_n47 <= '1';
   load_n_store_n46 <= '1';
   load_n_store_n45 <= '1';
   load_n_store_n44 <= '1';
   load_n_store_n43 <= '1';
   load_n_store_n42 <= '1';
   load_n_store_n41 <= '1';
   load_n_store_n40 <= '1';
   load_n_store_n39 <= '1';
   load_n_store_n38 <= '1';
   load_n_store_n37 <= '1';
   load_n_store_n36 <= '1';
   load_n_store_n35 <= '1';
   load_n_store_n34 <= '1';
   load_n_store_n33 <= '1';
   load_n_store_n32 <= '1';
   load_n_store_n31 <= '1';
   load_n_store_n30 <= '1';
   load_n_store_n29 <= '1';
   load_n_store_n28 <= '1';
   load_n_store_n27 <= '1';
   load_n_store_n26 <= '1';
   load_n_store_n25 <= '1';
   load_n_store_n24 <= '1';
   load_n_store_n23 <= '1';
   load_n_store_n22 <= '1';
   load_n_store_n21 <= '1';
   load_n_store_n20 <= '1';
   load_n_store_n19 <= '1';
   load_n_store_n18 <= '1';
   load_n_store_n17 <= '1';
   load_n_store_n16 <= '1';
   load_n_store_n15 <= '1';
   load_n_store_n14 <= '1';
   load_n_store_n13 <= '1';
   load_n_store_n12 <= '1';
   load_n_store_top_ack_reg : dff port map( d => load_n_store_n265, gclk => clk
                           , rnot => load_n_store_n12, q => top_ack_port);
   load_n_store_mem_out_b0_reg_7_inst : dff port map( d => n2241, gclk => clk, 
                           rnot => load_n_store_n13, q => mem_out_b0_7_port);
   load_n_store_mem_out_b0_reg_6_inst : dff port map( d => n2240, gclk => clk, 
                           rnot => load_n_store_n14, q => mem_out_b0_6_port);
   load_n_store_mem_out_b0_reg_5_inst : dff port map( d => n2239, gclk => clk, 
                           rnot => load_n_store_n15, q => mem_out_b0_5_port);
   load_n_store_mem_out_b0_reg_4_inst : dff port map( d => n2238, gclk => clk, 
                           rnot => load_n_store_n16, q => mem_out_b0_4_port);
   load_n_store_mem_out_b0_reg_3_inst : dff port map( d => n2237, gclk => clk, 
                           rnot => load_n_store_n17, q => mem_out_b0_3_port);
   load_n_store_mem_out_b0_reg_2_inst : dff port map( d => n2236, gclk => clk, 
                           rnot => load_n_store_n18, q => mem_out_b0_2_port);
   load_n_store_mem_out_b0_reg_1_inst : dff port map( d => n2235, gclk => clk, 
                           rnot => load_n_store_n19, q => mem_out_b0_1_port);
   load_n_store_mem_out_b0_reg_0_inst : dff port map( d => n2234, gclk => clk, 
                           rnot => load_n_store_n20, q => mem_out_b0_0_port);
   load_n_store_lazy_in_reg_0_7_inst : dff port map( d => n2265, gclk => clk, 
                           rnot => load_n_store_n21, q => 
                           load_n_store_lazy_in_0_7_port);
   load_n_store_lazy_in_reg_0_6_inst : dff port map( d => n2264, gclk => clk, 
                           rnot => load_n_store_n22, q => 
                           load_n_store_lazy_in_0_6_port);
   load_n_store_lazy_in_reg_0_5_inst : dff port map( d => n2263, gclk => clk, 
                           rnot => load_n_store_n23, q => 
                           load_n_store_lazy_in_0_5_port);
   load_n_store_lazy_in_reg_0_4_inst : dff port map( d => n2262, gclk => clk, 
                           rnot => load_n_store_n24, q => 
                           load_n_store_lazy_in_0_4_port);
   load_n_store_lazy_in_reg_0_3_inst : dff port map( d => n2261, gclk => clk, 
                           rnot => load_n_store_n25, q => 
                           load_n_store_lazy_in_0_3_port);
   load_n_store_lazy_in_reg_0_2_inst : dff port map( d => n2260, gclk => clk, 
                           rnot => load_n_store_n26, q => 
                           load_n_store_lazy_in_0_2_port);
   load_n_store_lazy_in_reg_0_1_inst : dff port map( d => n2259, gclk => clk, 
                           rnot => load_n_store_n27, q => 
                           load_n_store_lazy_in_0_1_port);
   load_n_store_lazy_in_reg_0_0_inst : dff port map( d => n2258, gclk => clk, 
                           rnot => load_n_store_n28, q => 
                           load_n_store_lazy_in_0_0_port);
   load_n_store_mem_out_g0_reg_7_inst : dff port map( d => n2233, gclk => clk, 
                           rnot => load_n_store_n29, q => mem_out_g0_7_port);
   load_n_store_mem_out_g0_reg_6_inst : dff port map( d => n2232, gclk => clk, 
                           rnot => load_n_store_n30, q => mem_out_g0_6_port);
   load_n_store_mem_out_g0_reg_5_inst : dff port map( d => n2231, gclk => clk, 
                           rnot => load_n_store_n31, q => mem_out_g0_5_port);
   load_n_store_mem_out_g0_reg_4_inst : dff port map( d => n2230, gclk => clk, 
                           rnot => load_n_store_n32, q => mem_out_g0_4_port);
   load_n_store_mem_out_g0_reg_3_inst : dff port map( d => n2229, gclk => clk, 
                           rnot => load_n_store_n33, q => mem_out_g0_3_port);
   load_n_store_mem_out_g0_reg_2_inst : dff port map( d => n2228, gclk => clk, 
                           rnot => load_n_store_n34, q => mem_out_g0_2_port);
   load_n_store_mem_out_g0_reg_1_inst : dff port map( d => n2227, gclk => clk, 
                           rnot => load_n_store_n35, q => mem_out_g0_1_port);
   load_n_store_mem_out_g0_reg_0_inst : dff port map( d => n2226, gclk => clk, 
                           rnot => load_n_store_n36, q => mem_out_g0_0_port);
   load_n_store_lazy_in_reg_1_7_inst : dff port map( d => n2257, gclk => clk, 
                           rnot => load_n_store_n37, q => 
                           load_n_store_lazy_in_1_7_port);
   load_n_store_lazy_in_reg_1_6_inst : dff port map( d => n2256, gclk => clk, 
                           rnot => load_n_store_n38, q => 
                           load_n_store_lazy_in_1_6_port);
   load_n_store_lazy_in_reg_1_5_inst : dff port map( d => n2255, gclk => clk, 
                           rnot => load_n_store_n39, q => 
                           load_n_store_lazy_in_1_5_port);
   load_n_store_lazy_in_reg_1_4_inst : dff port map( d => n2254, gclk => clk, 
                           rnot => load_n_store_n40, q => 
                           load_n_store_lazy_in_1_4_port);
   load_n_store_lazy_in_reg_1_3_inst : dff port map( d => n2253, gclk => clk, 
                           rnot => load_n_store_n41, q => 
                           load_n_store_lazy_in_1_3_port);
   load_n_store_lazy_in_reg_1_2_inst : dff port map( d => n2252, gclk => clk, 
                           rnot => load_n_store_n42, q => 
                           load_n_store_lazy_in_1_2_port);
   load_n_store_lazy_in_reg_1_1_inst : dff port map( d => n2251, gclk => clk, 
                           rnot => load_n_store_n43, q => 
                           load_n_store_lazy_in_1_1_port);
   load_n_store_lazy_in_reg_1_0_inst : dff port map( d => n2250, gclk => clk, 
                           rnot => load_n_store_n44, q => 
                           load_n_store_lazy_in_1_0_port);
   load_n_store_mem_out_r0_reg_7_inst : dff port map( d => n2225, gclk => clk, 
                           rnot => load_n_store_n45, q => mem_out_r0_7_port);
   load_n_store_mem_out_r0_reg_6_inst : dff port map( d => n2224, gclk => clk, 
                           rnot => load_n_store_n46, q => mem_out_r0_6_port);
   load_n_store_mem_out_r0_reg_5_inst : dff port map( d => n2223, gclk => clk, 
                           rnot => load_n_store_n47, q => mem_out_r0_5_port);
   load_n_store_mem_out_r0_reg_4_inst : dff port map( d => n2222, gclk => clk, 
                           rnot => load_n_store_n48, q => mem_out_r0_4_port);
   load_n_store_mem_out_r0_reg_3_inst : dff port map( d => n2221, gclk => clk, 
                           rnot => load_n_store_n49, q => mem_out_r0_3_port);
   load_n_store_mem_out_r0_reg_2_inst : dff port map( d => n2220, gclk => clk, 
                           rnot => load_n_store_n50, q => mem_out_r0_2_port);
   load_n_store_mem_out_r0_reg_1_inst : dff port map( d => n2219, gclk => clk, 
                           rnot => load_n_store_n51, q => mem_out_r0_1_port);
   load_n_store_mem_out_r0_reg_0_inst : dff port map( d => n2218, gclk => clk, 
                           rnot => load_n_store_n52, q => mem_out_r0_0_port);
   load_n_store_lazy_in_reg_2_7_inst : dff port map( d => n2249, gclk => clk, 
                           rnot => load_n_store_n53, q => 
                           load_n_store_lazy_in_2_7_port);
   load_n_store_lazy_in_reg_2_6_inst : dff port map( d => n2248, gclk => clk, 
                           rnot => load_n_store_n54, q => 
                           load_n_store_lazy_in_2_6_port);
   load_n_store_lazy_in_reg_2_5_inst : dff port map( d => n2247, gclk => clk, 
                           rnot => load_n_store_n55, q => 
                           load_n_store_lazy_in_2_5_port);
   load_n_store_lazy_in_reg_2_4_inst : dff port map( d => n2246, gclk => clk, 
                           rnot => load_n_store_n56, q => 
                           load_n_store_lazy_in_2_4_port);
   load_n_store_lazy_in_reg_2_3_inst : dff port map( d => n2245, gclk => clk, 
                           rnot => load_n_store_n57, q => 
                           load_n_store_lazy_in_2_3_port);
   load_n_store_lazy_in_reg_2_2_inst : dff port map( d => n2244, gclk => clk, 
                           rnot => load_n_store_n58, q => 
                           load_n_store_lazy_in_2_2_port);
   load_n_store_lazy_in_reg_2_1_inst : dff port map( d => n2243, gclk => clk, 
                           rnot => load_n_store_n59, q => 
                           load_n_store_lazy_in_2_1_port);
   load_n_store_lazy_in_reg_2_0_inst : dff port map( d => n2242, gclk => clk, 
                           rnot => load_n_store_n60, q => 
                           load_n_store_lazy_in_2_0_port);
   load_n_store_mem_reg_f_reg : dff port map( d => load_n_store_n259, gclk => 
                           clk, rnot => load_n_store_n61, q => mem_reg_f);
   load_n_store_mem_hub_f_reg : dff port map( d => load_n_store_n260, gclk => 
                           clk, rnot => load_n_store_n62, q => mem_hub_f);
   load_n_store_we_i_reg : dff port map( d => load_n_store_n264, gclk => clk, 
                           rnot => load_n_store_n63, q => load_n_store_we_i);
   load_n_store_simple_mem_sm_reg_1_inst : dff port map( d => load_n_store_n271
                           , gclk => clk, rnot => load_n_store_n64, q => 
                           load_n_store_simple_mem_sm_1_port);
   load_n_store_simple_mem_sm_reg_0_inst : dff port map( d => load_n_store_n266
                           , gclk => clk, rnot => load_n_store_n65, q => 
                           load_n_store_simple_mem_sm_0_port);
   load_n_store_mem_full_reg : dff port map( d => load_n_store_n272, gclk => 
                           clk, rnot => load_n_store_n66, q => 
                           load_n_store_mem_full);
   load_n_store_s_addr_reg_4_inst : dff port map( d => load_n_store_n273, gclk 
                           => clk, rnot => load_n_store_n67, q => 
                           load_n_store_s_addr_4_port);
   load_n_store_s_addr_reg_1_inst : dff port map( d => load_n_store_n263, gclk 
                           => clk, rnot => load_n_store_n68, q => 
                           load_n_store_s_addr_1_port);
   load_n_store_s_addr_reg_2_inst : dff port map( d => load_n_store_n262, gclk 
                           => clk, rnot => load_n_store_n69, q => 
                           load_n_store_s_addr_2_port);
   load_n_store_s_addr_reg_3_inst : dff port map( d => load_n_store_n261, gclk 
                           => clk, rnot => load_n_store_n70, q => 
                           load_n_store_s_addr_3_port);
   load_n_store_mem_timer_reg_0_inst : dff port map( d => load_n_store_n270, 
                           gclk => clk, rnot => load_n_store_n71, q => 
                           load_n_store_mem_timer_0_port);
   load_n_store_mem_timer_reg_1_inst : dff port map( d => load_n_store_n269, 
                           gclk => clk, rnot => load_n_store_n72, q => 
                           load_n_store_mem_timer_1_port);
   load_n_store_mem_timer_reg_2_inst : dff port map( d => load_n_store_n268, 
                           gclk => clk, rnot => load_n_store_n73, q => 
                           load_n_store_mem_timer_2_port);
   load_n_store_mem_timer_reg_3_inst : dff port map( d => load_n_store_n267, 
                           gclk => clk, rnot => load_n_store_n74, q => 
                           load_n_store_mem_timer_3_port);
   load_n_store_mem_timer_reg_4_inst : dff port map( d => load_n_store_n274, 
                           gclk => clk, rnot => load_n_store_n75, q => 
                           load_n_store_mem_timer_4_port);
   load_n_store_s_addr_reg_0_inst : dff port map( d => load_n_store_n275, gclk 
                           => clk, rnot => load_n_store_n76, q => 
                           load_n_store_s_addr_0_port);
   display_out_n151 <= '1';
   display_out_n150 <= '1';
   display_out_n149 <= '1';
   display_out_n148 <= '1';
   display_out_n147 <= '1';
   display_out_n146 <= '1';
   display_out_n145 <= '1';
   display_out_n144 <= '1';
   display_out_n143 <= '1';
   display_out_n142 <= '1';
   display_out_n141 <= '1';
   display_out_n140 <= '1';
   display_out_n139 <= '1';
   display_out_n138 <= '1';
   display_out_n137 <= '1';
   display_out_n136 <= '1';
   display_out_n135 <= '1';
   display_out_n134 <= '1';
   display_out_n133 <= '1';
   display_out_n132 <= '1';
   display_out_n131 <= '1';
   display_out_n130 <= '1';
   display_out_n129 <= '1';
   display_out_n128 <= '1';
   display_out_n127 <= '1';
   display_out_n126 <= '1';
   display_out_n125 <= '1';
   display_out_n124 <= '1';
   display_out_n123 <= '1';
   display_out_n122 <= '1';
   display_out_n121 <= '1';
   display_out_n120 <= '1';
   display_out_n119 <= '1';
   display_out_n118 <= '1';
   display_out_n117 <= '1';
   display_out_n116 <= '1';
   display_out_n115 <= '1';
   display_out_n114 <= '1';
   display_out_n113 <= '1';
   display_out_n112 <= '1';
   display_out_n111 <= '1';
   display_out_n110 <= '1';
   display_out_n109 <= '1';
   display_out_n108 <= '1';
   display_out_n107 <= '1';
   display_out_n106 <= '1';
   display_out_n105 <= '1';
   display_out_n104 <= '1';
   display_out_n103 <= '1';
   display_out_n102 <= '1';
   display_out_n101 <= '1';
   display_out_n100 <= '1';
   display_out_n99 <= '1';
   display_out_n98 <= '1';
   display_out_n97 <= '1';
   display_out_n96 <= '1';
   display_out_n95 <= '1';
   display_out_n94 <= '1';
   display_out_n93 <= '1';
   display_out_n92 <= '1';
   display_out_n91 <= '1';
   display_out_n90 <= '1';
   display_out_n89 <= '1';
   display_out_n88 <= '1';
   display_out_n87 <= '1';
   display_out_n86 <= '1';
   display_out_n85 <= '1';
   display_out_n84 <= '1';
   display_out_n83 <= '1';
   display_out_n82 <= '1';
   display_out_n81 <= '1';
   display_out_n80 <= '1';
   display_out_n79 <= '1';
   display_out_n78 <= '1';
   display_out_n77 <= '1';
   display_out_n76 <= '1';
   display_out_n75 <= '1';
   display_out_n74 <= '1';
   display_out_n73 <= '1';
   display_out_n72 <= '1';
   display_out_n71 <= '1';
   display_out_n70 <= '1';
   display_out_n69 <= '1';
   display_out_n68 <= '1';
   display_out_hub_b0_o_reg : dff port map( d => display_out_n474, gclk => clk,
                           rnot => display_out_n68, q => hub_b0_o_port);
   display_out_hub_g0_o_reg : dff port map( d => display_out_n475, gclk => clk,
                           rnot => display_out_n69, q => hub_g0_o_port);
   display_out_hub_r0_o_reg : dff port map( d => display_out_n476, gclk => clk,
                           rnot => display_out_n70, q => hub_r0_o_port);
   display_out_hub_piso_b0_reg_0_inst : dff port map( d => display_out_n477, 
                           gclk => clk, rnot => display_out_n71, q => 
                           display_out_hub_piso_b0_0_port);
   display_out_hub_piso_b0_reg_1_inst : dff port map( d => display_out_n483, 
                           gclk => clk, rnot => display_out_n72, q => 
                           display_out_hub_piso_b0_1_port);
   display_out_hub_piso_b0_reg_2_inst : dff port map( d => display_out_n482, 
                           gclk => clk, rnot => display_out_n73, q => 
                           display_out_hub_piso_b0_2_port);
   display_out_hub_piso_b0_reg_3_inst : dff port map( d => display_out_n481, 
                           gclk => clk, rnot => display_out_n74, q => 
                           display_out_hub_piso_b0_3_port);
   display_out_hub_piso_b0_reg_4_inst : dff port map( d => display_out_n480, 
                           gclk => clk, rnot => display_out_n75, q => 
                           display_out_hub_piso_b0_4_port);
   display_out_hub_piso_b0_reg_5_inst : dff port map( d => display_out_n479, 
                           gclk => clk, rnot => display_out_n76, q => 
                           display_out_hub_piso_b0_5_port);
   display_out_hub_piso_b0_reg_6_inst : dff port map( d => display_out_n478, 
                           gclk => clk, rnot => display_out_n77, q => 
                           display_out_hub_piso_b0_6_port);
   display_out_hub_piso_b0_reg_7_inst : dff port map( d => n2268, gclk => clk, 
                           rnot => display_out_n78, q => 
                           display_out_hub_piso_b0_7_port);
   display_out_hub_piso_g0_reg_0_inst : dff port map( d => display_out_n484, 
                           gclk => clk, rnot => display_out_n79, q => 
                           display_out_hub_piso_g0_0_port);
   display_out_hub_piso_g0_reg_1_inst : dff port map( d => display_out_n490, 
                           gclk => clk, rnot => display_out_n80, q => 
                           display_out_hub_piso_g0_1_port);
   display_out_hub_piso_g0_reg_2_inst : dff port map( d => display_out_n489, 
                           gclk => clk, rnot => display_out_n81, q => 
                           display_out_hub_piso_g0_2_port);
   display_out_hub_piso_g0_reg_3_inst : dff port map( d => display_out_n488, 
                           gclk => clk, rnot => display_out_n82, q => 
                           display_out_hub_piso_g0_3_port);
   display_out_hub_piso_g0_reg_4_inst : dff port map( d => display_out_n487, 
                           gclk => clk, rnot => display_out_n83, q => 
                           display_out_hub_piso_g0_4_port);
   display_out_hub_piso_g0_reg_5_inst : dff port map( d => display_out_n486, 
                           gclk => clk, rnot => display_out_n84, q => 
                           display_out_hub_piso_g0_5_port);
   display_out_hub_piso_g0_reg_6_inst : dff port map( d => display_out_n485, 
                           gclk => clk, rnot => display_out_n85, q => 
                           display_out_hub_piso_g0_6_port);
   display_out_hub_piso_g0_reg_7_inst : dff port map( d => n2266, gclk => clk, 
                           rnot => display_out_n86, q => 
                           display_out_hub_piso_g0_7_port);
   display_out_hub_piso_r0_reg_0_inst : dff port map( d => display_out_n491, 
                           gclk => clk, rnot => display_out_n87, q => 
                           display_out_hub_piso_r0_0_port);
   display_out_hub_piso_r0_reg_1_inst : dff port map( d => display_out_n497, 
                           gclk => clk, rnot => display_out_n88, q => 
                           display_out_hub_piso_r0_1_port);
   display_out_hub_piso_r0_reg_2_inst : dff port map( d => display_out_n496, 
                           gclk => clk, rnot => display_out_n89, q => 
                           display_out_hub_piso_r0_2_port);
   display_out_hub_piso_r0_reg_3_inst : dff port map( d => display_out_n495, 
                           gclk => clk, rnot => display_out_n90, q => 
                           display_out_hub_piso_r0_3_port);
   display_out_hub_piso_r0_reg_4_inst : dff port map( d => display_out_n494, 
                           gclk => clk, rnot => display_out_n91, q => 
                           display_out_hub_piso_r0_4_port);
   display_out_hub_piso_r0_reg_5_inst : dff port map( d => display_out_n493, 
                           gclk => clk, rnot => display_out_n92, q => 
                           display_out_hub_piso_r0_5_port);
   display_out_hub_piso_r0_reg_6_inst : dff port map( d => display_out_n492, 
                           gclk => clk, rnot => display_out_n93, q => 
                           display_out_hub_piso_r0_6_port);
   display_out_hub_piso_r0_reg_7_inst : dff port map( d => n2267, gclk => clk, 
                           rnot => display_out_n94, q => 
                           display_out_hub_piso_r0_7_port);
   display_out_hub_blank_o_reg : dff port map( d => display_out_n508, gclk => 
                           clk, rnot => display_out_n95, q => hub_blank_o_port)
                           ;
   display_out_hub_mux_o_reg_1_inst : dff port map( d => display_out_n503, gclk
                           => clk, rnot => display_out_n96, q => 
                           hub_mux_o_1_port);
   display_out_hub_mux_o_reg_0_inst : dff port map( d => display_out_n504, gclk
                           => clk, rnot => display_out_n97, q => 
                           hub_mux_o_0_port);
   display_out_hub_mux_o_reg_2_inst : dff port map( d => display_out_n507, gclk
                           => clk, rnot => display_out_n98, q => 
                           hub_mux_o_2_port);
   display_out_h_row_reg_1_inst : dff port map( d => display_out_n505, gclk => 
                           clk, rnot => display_out_n99, q => 
                           display_out_h_row_1_port);
   display_out_h_row_reg_0_inst : dff port map( d => display_out_n506, gclk => 
                           clk, rnot => display_out_n100, q => 
                           display_out_h_row_0_port);
   display_out_hub_latch_o_reg : dff port map( d => display_out_n498, gclk => 
                           clk, rnot => display_out_n101, q => hub_latch_o_port
                           );
   display_out_hub_clk_o_reg : dff port map( d => display_out_n502, gclk => clk
                           , rnot => display_out_n102, q => hub_clk_o_port);
   display_out_hub_reg_f_reg : dff port map( d => display_out_n501, gclk => clk
                           , rnot => display_out_n103, q => hub_reg_f);
   display_out_disp_timer_reg_31_inst : dff port map( d => n2273, gclk => clk, 
                           rnot => display_out_n104, q => 
                           display_out_disp_timer_31_port);
   display_out_disp_timer_reg_30_inst : dff port map( d => n2274, gclk => clk, 
                           rnot => display_out_n105, q => 
                           display_out_disp_timer_30_port);
   display_out_disp_timer_reg_29_inst : dff port map( d => n2275, gclk => clk, 
                           rnot => display_out_n106, q => 
                           display_out_disp_timer_29_port);
   display_out_disp_timer_reg_28_inst : dff port map( d => n2276, gclk => clk, 
                           rnot => display_out_n107, q => 
                           display_out_disp_timer_28_port);
   display_out_disp_timer_reg_27_inst : dff port map( d => n2277, gclk => clk, 
                           rnot => display_out_n108, q => 
                           display_out_disp_timer_27_port);
   display_out_disp_timer_reg_26_inst : dff port map( d => n2278, gclk => clk, 
                           rnot => display_out_n109, q => 
                           display_out_disp_timer_26_port);
   display_out_disp_timer_reg_25_inst : dff port map( d => n2279, gclk => clk, 
                           rnot => display_out_n110, q => 
                           display_out_disp_timer_25_port);
   display_out_disp_timer_reg_24_inst : dff port map( d => n2280, gclk => clk, 
                           rnot => display_out_n111, q => 
                           display_out_disp_timer_24_port);
   display_out_disp_timer_reg_23_inst : dff port map( d => n2281, gclk => clk, 
                           rnot => display_out_n112, q => 
                           display_out_disp_timer_23_port);
   display_out_disp_timer_reg_22_inst : dff port map( d => n2282, gclk => clk, 
                           rnot => display_out_n113, q => 
                           display_out_disp_timer_22_port);
   display_out_disp_timer_reg_21_inst : dff port map( d => n2283, gclk => clk, 
                           rnot => display_out_n114, q => 
                           display_out_disp_timer_21_port);
   display_out_disp_timer_reg_20_inst : dff port map( d => n2284, gclk => clk, 
                           rnot => display_out_n115, q => 
                           display_out_disp_timer_20_port);
   display_out_disp_timer_reg_19_inst : dff port map( d => n2285, gclk => clk, 
                           rnot => display_out_n116, q => 
                           display_out_disp_timer_19_port);
   display_out_disp_timer_reg_18_inst : dff port map( d => n2286, gclk => clk, 
                           rnot => display_out_n117, q => 
                           display_out_disp_timer_18_port);
   display_out_disp_timer_reg_17_inst : dff port map( d => n2287, gclk => clk, 
                           rnot => display_out_n118, q => 
                           display_out_disp_timer_17_port);
   display_out_disp_timer_reg_16_inst : dff port map( d => n2288, gclk => clk, 
                           rnot => display_out_n119, q => 
                           display_out_disp_timer_16_port);
   display_out_disp_timer_reg_15_inst : dff port map( d => display_out_n525, 
                           gclk => clk, rnot => display_out_n120, q => 
                           display_out_disp_timer_15_port);
   display_out_disp_timer_reg_14_inst : dff port map( d => display_out_n524, 
                           gclk => clk, rnot => display_out_n121, q => 
                           display_out_disp_timer_14_port);
   display_out_disp_timer_reg_13_inst : dff port map( d => display_out_n523, 
                           gclk => clk, rnot => display_out_n122, q => 
                           display_out_disp_timer_13_port);
   display_out_disp_timer_reg_12_inst : dff port map( d => display_out_n522, 
                           gclk => clk, rnot => display_out_n123, q => 
                           display_out_disp_timer_12_port);
   display_out_disp_timer_reg_11_inst : dff port map( d => display_out_n521, 
                           gclk => clk, rnot => display_out_n124, q => 
                           display_out_disp_timer_11_port);
   display_out_disp_timer_reg_10_inst : dff port map( d => display_out_n520, 
                           gclk => clk, rnot => display_out_n125, q => 
                           display_out_disp_timer_10_port);
   display_out_disp_timer_reg_9_inst : dff port map( d => display_out_n519, 
                           gclk => clk, rnot => display_out_n126, q => 
                           display_out_disp_timer_9_port);
   display_out_disp_timer_reg_7_inst : dff port map( d => display_out_n517, 
                           gclk => clk, rnot => display_out_n127, q => 
                           display_out_disp_timer_7_port);
   display_out_disp_timer_reg_6_inst : dff port map( d => display_out_n516, 
                           gclk => clk, rnot => display_out_n128, q => 
                           display_out_disp_timer_6_port);
   display_out_disp_timer_reg_5_inst : dff port map( d => display_out_n515, 
                           gclk => clk, rnot => display_out_n129, q => 
                           display_out_disp_timer_5_port);
   display_out_disp_timer_reg_3_inst : dff port map( d => display_out_n513, 
                           gclk => clk, rnot => display_out_n130, q => 
                           display_out_disp_timer_3_port);
   display_out_disp_timer_reg_1_inst : dff port map( d => display_out_n511, 
                           gclk => clk, rnot => display_out_n131, q => 
                           display_out_disp_timer_1_port);
   display_out_disp_timer_reg_0_inst : dff port map( d => display_out_n526, 
                           gclk => clk, rnot => display_out_n132, q => 
                           display_out_disp_timer_0_port);
   display_out_disp_timer_reg_8_inst : dff port map( d => display_out_n518, 
                           gclk => clk, rnot => display_out_n133, q => 
                           display_out_disp_timer_8_port);
   display_out_bcd_time_reg_1_inst : dff port map( d => display_out_n509, gclk 
                           => clk, rnot => display_out_n134, q => 
                           display_out_bcd_time_1_port);
   display_out_h_col_reg_1_inst : dff port map( d => display_out_n533, gclk => 
                           clk, rnot => display_out_n135, q => 
                           display_out_h_col_1_port);
   display_out_bcd_time_reg_0_inst : dff port map( d => display_out_n510, gclk 
                           => clk, rnot => display_out_n136, q => 
                           display_out_bcd_time_0_port);
   display_out_h_col_reg_0_inst : dff port map( d => display_out_n500, gclk => 
                           clk, rnot => display_out_n137, q => 
                           display_out_h_col_0_port);
   display_out_clk_timer_reg_6_inst : dff port map( d => n2269, gclk => clk, 
                           rnot => display_out_n138, q => 
                           display_out_clk_timer_6_port);
   display_out_clk_timer_reg_5_inst : dff port map( d => n2270, gclk => clk, 
                           rnot => display_out_n139, q => 
                           display_out_clk_timer_5_port);
   display_out_clk_timer_reg_4_inst : dff port map( d => display_out_n529, gclk
                           => clk, rnot => display_out_n140, q => 
                           display_out_clk_timer_4_port);
   display_out_clk_timer_reg_3_inst : dff port map( d => display_out_n528, gclk
                           => clk, rnot => display_out_n141, q => 
                           display_out_clk_timer_3_port);
   display_out_clk_timer_reg_2_inst : dff port map( d => display_out_n527, gclk
                           => clk, rnot => display_out_n142, q => 
                           display_out_clk_timer_2_port);
   display_out_clk_timer_reg_1_inst : dff port map( d => n2271, gclk => clk, 
                           rnot => display_out_n143, q => 
                           display_out_clk_timer_1_port);
   display_out_clk_timer_reg_0_inst : dff port map( d => display_out_n530, gclk
                           => clk, rnot => display_out_n144, q => 
                           display_out_clk_timer_0_port);
   display_out_h_col_reg_2_inst : dff port map( d => display_out_n499, gclk => 
                           clk, rnot => display_out_n145, q => 
                           display_out_h_col_2_port);
   display_out_disp_timer_reg_2_inst : dff port map( d => display_out_n512, 
                           gclk => clk, rnot => display_out_n146, q => 
                           display_out_disp_timer_2_port);
   display_out_bcd_time_reg_2_inst : dff port map( d => display_out_n532, gclk 
                           => clk, rnot => display_out_n147, q => 
                           display_out_bcd_time_2_port);
   display_out_hub_out_sm_reg_2_inst : dff port map( d => display_out_n534, 
                           gclk => clk, rnot => display_out_n148, q => 
                           display_out_hub_out_sm_2_port);
   display_out_disp_timer_reg_4_inst : dff port map( d => display_out_n514, 
                           gclk => clk, rnot => display_out_n149, q => 
                           display_out_disp_timer_4_port);
   display_out_hub_out_sm_reg_1_inst : dff port map( d => display_out_n531, 
                           gclk => clk, rnot => display_out_n150, q => 
                           display_out_hub_out_sm_1_port);
   display_out_hub_out_sm_reg_0_inst : dff port map( d => display_out_n535, 
                           gclk => clk, rnot => display_out_n151, q => 
                           display_out_hub_out_sm_0_port);
   load_n_store_RGB_Array_0_n906 <= '1';
   load_n_store_RGB_Array_0_n905 <= '1';
   load_n_store_RGB_Array_0_n904 <= '1';
   load_n_store_RGB_Array_0_n903 <= '1';
   load_n_store_RGB_Array_0_n902 <= '1';
   load_n_store_RGB_Array_0_n901 <= '1';
   load_n_store_RGB_Array_0_n900 <= '1';
   load_n_store_RGB_Array_0_n899 <= '1';
   load_n_store_RGB_Array_0_n898 <= '1';
   load_n_store_RGB_Array_0_n897 <= '1';
   load_n_store_RGB_Array_0_n896 <= '1';
   load_n_store_RGB_Array_0_n895 <= '1';
   load_n_store_RGB_Array_0_n894 <= '1';
   load_n_store_RGB_Array_0_n893 <= '1';
   load_n_store_RGB_Array_0_n892 <= '1';
   load_n_store_RGB_Array_0_n891 <= '1';
   load_n_store_RGB_Array_0_n890 <= '1';
   load_n_store_RGB_Array_0_n889 <= '1';
   load_n_store_RGB_Array_0_n888 <= '1';
   load_n_store_RGB_Array_0_n887 <= '1';
   load_n_store_RGB_Array_0_n886 <= '1';
   load_n_store_RGB_Array_0_n885 <= '1';
   load_n_store_RGB_Array_0_n884 <= '1';
   load_n_store_RGB_Array_0_n883 <= '1';
   load_n_store_RGB_Array_0_n882 <= '1';
   load_n_store_RGB_Array_0_n881 <= '1';
   load_n_store_RGB_Array_0_n880 <= '1';
   load_n_store_RGB_Array_0_n879 <= '1';
   load_n_store_RGB_Array_0_n878 <= '1';
   load_n_store_RGB_Array_0_n877 <= '1';
   load_n_store_RGB_Array_0_n876 <= '1';
   load_n_store_RGB_Array_0_n875 <= '1';
   load_n_store_RGB_Array_0_n874 <= '1';
   load_n_store_RGB_Array_0_n873 <= '1';
   load_n_store_RGB_Array_0_n872 <= '1';
   load_n_store_RGB_Array_0_n871 <= '1';
   load_n_store_RGB_Array_0_n870 <= '1';
   load_n_store_RGB_Array_0_n869 <= '1';
   load_n_store_RGB_Array_0_n868 <= '1';
   load_n_store_RGB_Array_0_n867 <= '1';
   load_n_store_RGB_Array_0_n866 <= '1';
   load_n_store_RGB_Array_0_n865 <= '1';
   load_n_store_RGB_Array_0_n864 <= '1';
   load_n_store_RGB_Array_0_n863 <= '1';
   load_n_store_RGB_Array_0_n862 <= '1';
   load_n_store_RGB_Array_0_n861 <= '1';
   load_n_store_RGB_Array_0_n860 <= '1';
   load_n_store_RGB_Array_0_n859 <= '1';
   load_n_store_RGB_Array_0_n858 <= '1';
   load_n_store_RGB_Array_0_n857 <= '1';
   load_n_store_RGB_Array_0_n856 <= '1';
   load_n_store_RGB_Array_0_n855 <= '1';
   load_n_store_RGB_Array_0_n854 <= '1';
   load_n_store_RGB_Array_0_n853 <= '1';
   load_n_store_RGB_Array_0_n852 <= '1';
   load_n_store_RGB_Array_0_n851 <= '1';
   load_n_store_RGB_Array_0_n850 <= '1';
   load_n_store_RGB_Array_0_n849 <= '1';
   load_n_store_RGB_Array_0_n848 <= '1';
   load_n_store_RGB_Array_0_n847 <= '1';
   load_n_store_RGB_Array_0_n846 <= '1';
   load_n_store_RGB_Array_0_n845 <= '1';
   load_n_store_RGB_Array_0_n844 <= '1';
   load_n_store_RGB_Array_0_n843 <= '1';
   load_n_store_RGB_Array_0_n842 <= '1';
   load_n_store_RGB_Array_0_n841 <= '1';
   load_n_store_RGB_Array_0_n840 <= '1';
   load_n_store_RGB_Array_0_n839 <= '1';
   load_n_store_RGB_Array_0_n838 <= '1';
   load_n_store_RGB_Array_0_n837 <= '1';
   load_n_store_RGB_Array_0_n836 <= '1';
   load_n_store_RGB_Array_0_n835 <= '1';
   load_n_store_RGB_Array_0_n834 <= '1';
   load_n_store_RGB_Array_0_n833 <= '1';
   load_n_store_RGB_Array_0_n832 <= '1';
   load_n_store_RGB_Array_0_n831 <= '1';
   load_n_store_RGB_Array_0_n830 <= '1';
   load_n_store_RGB_Array_0_n829 <= '1';
   load_n_store_RGB_Array_0_n828 <= '1';
   load_n_store_RGB_Array_0_n827 <= '1';
   load_n_store_RGB_Array_0_n826 <= '1';
   load_n_store_RGB_Array_0_n825 <= '1';
   load_n_store_RGB_Array_0_n824 <= '1';
   load_n_store_RGB_Array_0_n823 <= '1';
   load_n_store_RGB_Array_0_n822 <= '1';
   load_n_store_RGB_Array_0_n821 <= '1';
   load_n_store_RGB_Array_0_n820 <= '1';
   load_n_store_RGB_Array_0_n819 <= '1';
   load_n_store_RGB_Array_0_n818 <= '1';
   load_n_store_RGB_Array_0_n817 <= '1';
   load_n_store_RGB_Array_0_n816 <= '1';
   load_n_store_RGB_Array_0_n815 <= '1';
   load_n_store_RGB_Array_0_n814 <= '1';
   load_n_store_RGB_Array_0_n813 <= '1';
   load_n_store_RGB_Array_0_n812 <= '1';
   load_n_store_RGB_Array_0_n811 <= '1';
   load_n_store_RGB_Array_0_n810 <= '1';
   load_n_store_RGB_Array_0_n809 <= '1';
   load_n_store_RGB_Array_0_n808 <= '1';
   load_n_store_RGB_Array_0_n807 <= '1';
   load_n_store_RGB_Array_0_n806 <= '1';
   load_n_store_RGB_Array_0_n805 <= '1';
   load_n_store_RGB_Array_0_n804 <= '1';
   load_n_store_RGB_Array_0_n803 <= '1';
   load_n_store_RGB_Array_0_n802 <= '1';
   load_n_store_RGB_Array_0_n801 <= '1';
   load_n_store_RGB_Array_0_n800 <= '1';
   load_n_store_RGB_Array_0_n799 <= '1';
   load_n_store_RGB_Array_0_n798 <= '1';
   load_n_store_RGB_Array_0_n797 <= '1';
   load_n_store_RGB_Array_0_n796 <= '1';
   load_n_store_RGB_Array_0_n795 <= '1';
   load_n_store_RGB_Array_0_n794 <= '1';
   load_n_store_RGB_Array_0_n793 <= '1';
   load_n_store_RGB_Array_0_n792 <= '1';
   load_n_store_RGB_Array_0_n791 <= '1';
   load_n_store_RGB_Array_0_n790 <= '1';
   load_n_store_RGB_Array_0_n789 <= '1';
   load_n_store_RGB_Array_0_n788 <= '1';
   load_n_store_RGB_Array_0_n787 <= '1';
   load_n_store_RGB_Array_0_n786 <= '1';
   load_n_store_RGB_Array_0_n785 <= '1';
   load_n_store_RGB_Array_0_n784 <= '1';
   load_n_store_RGB_Array_0_n783 <= '1';
   load_n_store_RGB_Array_0_n782 <= '1';
   load_n_store_RGB_Array_0_n781 <= '1';
   load_n_store_RGB_Array_0_n780 <= '1';
   load_n_store_RGB_Array_0_n779 <= '1';
   load_n_store_RGB_Array_0_n778 <= '1';
   load_n_store_RGB_Array_0_n777 <= '1';
   load_n_store_RGB_Array_0_n776 <= '1';
   load_n_store_RGB_Array_0_n775 <= '1';
   load_n_store_RGB_Array_0_n774 <= '1';
   load_n_store_RGB_Array_0_n773 <= '1';
   load_n_store_RGB_Array_0_n772 <= '1';
   load_n_store_RGB_Array_0_n771 <= '1';
   load_n_store_RGB_Array_0_n770 <= '1';
   load_n_store_RGB_Array_0_n769 <= '1';
   load_n_store_RGB_Array_0_n768 <= '1';
   load_n_store_RGB_Array_0_n767 <= '1';
   load_n_store_RGB_Array_0_n766 <= '1';
   load_n_store_RGB_Array_0_n765 <= '1';
   load_n_store_RGB_Array_0_n764 <= '1';
   load_n_store_RGB_Array_0_n763 <= '1';
   load_n_store_RGB_Array_0_n762 <= '1';
   load_n_store_RGB_Array_0_n761 <= '1';
   load_n_store_RGB_Array_0_n760 <= '1';
   load_n_store_RGB_Array_0_n759 <= '1';
   load_n_store_RGB_Array_0_n758 <= '1';
   load_n_store_RGB_Array_0_n757 <= '1';
   load_n_store_RGB_Array_0_n756 <= '1';
   load_n_store_RGB_Array_0_n755 <= '1';
   load_n_store_RGB_Array_0_n754 <= '1';
   load_n_store_RGB_Array_0_n753 <= '1';
   load_n_store_RGB_Array_0_n752 <= '1';
   load_n_store_RGB_Array_0_n751 <= '1';
   load_n_store_RGB_Array_0_n750 <= '1';
   load_n_store_RGB_Array_0_n749 <= '1';
   load_n_store_RGB_Array_0_n748 <= '1';
   load_n_store_RGB_Array_0_n747 <= '1';
   load_n_store_RGB_Array_0_n746 <= '1';
   load_n_store_RGB_Array_0_n745 <= '1';
   load_n_store_RGB_Array_0_n744 <= '1';
   load_n_store_RGB_Array_0_n743 <= '1';
   load_n_store_RGB_Array_0_n742 <= '1';
   load_n_store_RGB_Array_0_n741 <= '1';
   load_n_store_RGB_Array_0_n740 <= '1';
   load_n_store_RGB_Array_0_n739 <= '1';
   load_n_store_RGB_Array_0_n738 <= '1';
   load_n_store_RGB_Array_0_n737 <= '1';
   load_n_store_RGB_Array_0_n736 <= '1';
   load_n_store_RGB_Array_0_n735 <= '1';
   load_n_store_RGB_Array_0_n734 <= '1';
   load_n_store_RGB_Array_0_n733 <= '1';
   load_n_store_RGB_Array_0_n732 <= '1';
   load_n_store_RGB_Array_0_n731 <= '1';
   load_n_store_RGB_Array_0_n730 <= '1';
   load_n_store_RGB_Array_0_n729 <= '1';
   load_n_store_RGB_Array_0_n728 <= '1';
   load_n_store_RGB_Array_0_n727 <= '1';
   load_n_store_RGB_Array_0_n726 <= '1';
   load_n_store_RGB_Array_0_n725 <= '1';
   load_n_store_RGB_Array_0_n724 <= '1';
   load_n_store_RGB_Array_0_n723 <= '1';
   load_n_store_RGB_Array_0_n722 <= '1';
   load_n_store_RGB_Array_0_n721 <= '1';
   load_n_store_RGB_Array_0_n720 <= '1';
   load_n_store_RGB_Array_0_n719 <= '1';
   load_n_store_RGB_Array_0_n718 <= '1';
   load_n_store_RGB_Array_0_n717 <= '1';
   load_n_store_RGB_Array_0_n716 <= '1';
   load_n_store_RGB_Array_0_n715 <= '1';
   load_n_store_RGB_Array_0_n714 <= '1';
   load_n_store_RGB_Array_0_n713 <= '1';
   load_n_store_RGB_Array_0_n712 <= '1';
   load_n_store_RGB_Array_0_n711 <= '1';
   load_n_store_RGB_Array_0_n710 <= '1';
   load_n_store_RGB_Array_0_n709 <= '1';
   load_n_store_RGB_Array_0_n708 <= '1';
   load_n_store_RGB_Array_0_n707 <= '1';
   load_n_store_RGB_Array_0_n706 <= '1';
   load_n_store_RGB_Array_0_n705 <= '1';
   load_n_store_RGB_Array_0_n704 <= '1';
   load_n_store_RGB_Array_0_n703 <= '1';
   load_n_store_RGB_Array_0_n702 <= '1';
   load_n_store_RGB_Array_0_n701 <= '1';
   load_n_store_RGB_Array_0_n700 <= '1';
   load_n_store_RGB_Array_0_n699 <= '1';
   load_n_store_RGB_Array_0_n698 <= '1';
   load_n_store_RGB_Array_0_n697 <= '1';
   load_n_store_RGB_Array_0_n696 <= '1';
   load_n_store_RGB_Array_0_n695 <= '1';
   load_n_store_RGB_Array_0_n694 <= '1';
   load_n_store_RGB_Array_0_n693 <= '1';
   load_n_store_RGB_Array_0_n692 <= '1';
   load_n_store_RGB_Array_0_n691 <= '1';
   load_n_store_RGB_Array_0_n690 <= '1';
   load_n_store_RGB_Array_0_n689 <= '1';
   load_n_store_RGB_Array_0_n688 <= '1';
   load_n_store_RGB_Array_0_n687 <= '1';
   load_n_store_RGB_Array_0_n686 <= '1';
   load_n_store_RGB_Array_0_n685 <= '1';
   load_n_store_RGB_Array_0_n684 <= '1';
   load_n_store_RGB_Array_0_n683 <= '1';
   load_n_store_RGB_Array_0_n682 <= '1';
   load_n_store_RGB_Array_0_n681 <= '1';
   load_n_store_RGB_Array_0_n680 <= '1';
   load_n_store_RGB_Array_0_n679 <= '1';
   load_n_store_RGB_Array_0_n678 <= '1';
   load_n_store_RGB_Array_0_n677 <= '1';
   load_n_store_RGB_Array_0_n676 <= '1';
   load_n_store_RGB_Array_0_n675 <= '1';
   load_n_store_RGB_Array_0_n674 <= '1';
   load_n_store_RGB_Array_0_n673 <= '1';
   load_n_store_RGB_Array_0_n672 <= '1';
   load_n_store_RGB_Array_0_n671 <= '1';
   load_n_store_RGB_Array_0_n670 <= '1';
   load_n_store_RGB_Array_0_n669 <= '1';
   load_n_store_RGB_Array_0_n668 <= '1';
   load_n_store_RGB_Array_0_n667 <= '1';
   load_n_store_RGB_Array_0_n666 <= '1';
   load_n_store_RGB_Array_0_n665 <= '1';
   load_n_store_RGB_Array_0_n664 <= '1';
   load_n_store_RGB_Array_0_n663 <= '1';
   load_n_store_RGB_Array_0_n662 <= '1';
   load_n_store_RGB_Array_0_n661 <= '1';
   load_n_store_RGB_Array_0_n660 <= '1';
   load_n_store_RGB_Array_0_n659 <= '1';
   load_n_store_RGB_Array_0_n658 <= '1';
   load_n_store_RGB_Array_0_n656 <= '1';
   load_n_store_RGB_Array_0_n655 <= '1';
   load_n_store_RGB_Array_0_n653 <= '1';
   load_n_store_RGB_Array_0_n652 <= '1';
   load_n_store_RGB_Array_0_n650 <= '1';
   load_n_store_RGB_Array_0_n649 <= '1';
   load_n_store_RGB_Array_0_n647 <= '1';
   load_n_store_RGB_Array_0_n646 <= '1';
   load_n_store_RGB_Array_0_n644 <= '1';
   load_n_store_RGB_Array_0_n643 <= '1';
   load_n_store_RGB_Array_0_n641 <= '1';
   load_n_store_RGB_Array_0_n640 <= '1';
   load_n_store_RGB_Array_0_n638 <= '1';
   load_n_store_RGB_Array_0_n637 <= '1';
   load_n_store_RGB_Array_0_n635 <= '1';
   load_n_store_RGB_Array_0_data_out_o_reg_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n636, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n635, q => 
                           load_n_store_lazy_out_0_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_0_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n907, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n637, q => 
                           load_n_store_RGB_Array_0_block_ram_r_0_0_port);
   load_n_store_RGB_Array_0_data_out_o_reg_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n639, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n638, q => 
                           load_n_store_lazy_out_0_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_0_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n908, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n640, q => 
                           load_n_store_RGB_Array_0_block_ram_r_0_1_port);
   load_n_store_RGB_Array_0_data_out_o_reg_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n642, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n641, q => 
                           load_n_store_lazy_out_0_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_0_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n909, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n643, q => 
                           load_n_store_RGB_Array_0_block_ram_r_0_2_port);
   load_n_store_RGB_Array_0_data_out_o_reg_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n645, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n644, q => 
                           load_n_store_lazy_out_0_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_0_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n910, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n646, q => 
                           load_n_store_RGB_Array_0_block_ram_r_0_3_port);
   load_n_store_RGB_Array_0_data_out_o_reg_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n648, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n647, q => 
                           load_n_store_lazy_out_0_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_0_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n911, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n649, q => 
                           load_n_store_RGB_Array_0_block_ram_r_0_4_port);
   load_n_store_RGB_Array_0_data_out_o_reg_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n651, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n650, q => 
                           load_n_store_lazy_out_0_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_0_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n912, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n652, q => 
                           load_n_store_RGB_Array_0_block_ram_r_0_5_port);
   load_n_store_RGB_Array_0_data_out_o_reg_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n654, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n653, q => 
                           load_n_store_lazy_out_0_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_0_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n913, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n655, q => 
                           load_n_store_RGB_Array_0_block_ram_r_0_6_port);
   load_n_store_RGB_Array_0_data_out_o_reg_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n657, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n656, q => 
                           load_n_store_lazy_out_0_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_0_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n914, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n658, q => 
                           load_n_store_RGB_Array_0_block_ram_r_0_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_1_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n915, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n659, q => 
                           load_n_store_RGB_Array_0_block_ram_r_1_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_1_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n916, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n660, q => 
                           load_n_store_RGB_Array_0_block_ram_r_1_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_1_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n917, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n661, q => 
                           load_n_store_RGB_Array_0_block_ram_r_1_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_1_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n918, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n662, q => 
                           load_n_store_RGB_Array_0_block_ram_r_1_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_1_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n919, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n663, q => 
                           load_n_store_RGB_Array_0_block_ram_r_1_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_1_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n920, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n664, q => 
                           load_n_store_RGB_Array_0_block_ram_r_1_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_1_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n921, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n665, q => 
                           load_n_store_RGB_Array_0_block_ram_r_1_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_1_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n922, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n666, q => 
                           load_n_store_RGB_Array_0_block_ram_r_1_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_2_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n923, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n667, q => 
                           load_n_store_RGB_Array_0_block_ram_r_2_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_2_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n924, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n668, q => 
                           load_n_store_RGB_Array_0_block_ram_r_2_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_2_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n925, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n669, q => 
                           load_n_store_RGB_Array_0_block_ram_r_2_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_2_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n926, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n670, q => 
                           load_n_store_RGB_Array_0_block_ram_r_2_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_2_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n927, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n671, q => 
                           load_n_store_RGB_Array_0_block_ram_r_2_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_2_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n928, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n672, q => 
                           load_n_store_RGB_Array_0_block_ram_r_2_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_2_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n929, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n673, q => 
                           load_n_store_RGB_Array_0_block_ram_r_2_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_2_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n930, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n674, q => 
                           load_n_store_RGB_Array_0_block_ram_r_2_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_3_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n931, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n675, q => 
                           load_n_store_RGB_Array_0_block_ram_r_3_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_3_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n932, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n676, q => 
                           load_n_store_RGB_Array_0_block_ram_r_3_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_3_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n933, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n677, q => 
                           load_n_store_RGB_Array_0_block_ram_r_3_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_3_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n934, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n678, q => 
                           load_n_store_RGB_Array_0_block_ram_r_3_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_3_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n935, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n679, q => 
                           load_n_store_RGB_Array_0_block_ram_r_3_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_3_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n936, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n680, q => 
                           load_n_store_RGB_Array_0_block_ram_r_3_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_3_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n937, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n681, q => 
                           load_n_store_RGB_Array_0_block_ram_r_3_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_3_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n938, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n682, q => 
                           load_n_store_RGB_Array_0_block_ram_r_3_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_4_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n939, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n683, q => 
                           load_n_store_RGB_Array_0_block_ram_r_4_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_4_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n940, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n684, q => 
                           load_n_store_RGB_Array_0_block_ram_r_4_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_4_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n941, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n685, q => 
                           load_n_store_RGB_Array_0_block_ram_r_4_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_4_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n942, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n686, q => 
                           load_n_store_RGB_Array_0_block_ram_r_4_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_4_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n943, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n687, q => 
                           load_n_store_RGB_Array_0_block_ram_r_4_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_4_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n944, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n688, q => 
                           load_n_store_RGB_Array_0_block_ram_r_4_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_4_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n945, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n689, q => 
                           load_n_store_RGB_Array_0_block_ram_r_4_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_4_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n946, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n690, q => 
                           load_n_store_RGB_Array_0_block_ram_r_4_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_5_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n947, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n691, q => 
                           load_n_store_RGB_Array_0_block_ram_r_5_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_5_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n948, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n692, q => 
                           load_n_store_RGB_Array_0_block_ram_r_5_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_5_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n949, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n693, q => 
                           load_n_store_RGB_Array_0_block_ram_r_5_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_5_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n950, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n694, q => 
                           load_n_store_RGB_Array_0_block_ram_r_5_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_5_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n951, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n695, q => 
                           load_n_store_RGB_Array_0_block_ram_r_5_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_5_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n952, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n696, q => 
                           load_n_store_RGB_Array_0_block_ram_r_5_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_5_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n953, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n697, q => 
                           load_n_store_RGB_Array_0_block_ram_r_5_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_5_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n954, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n698, q => 
                           load_n_store_RGB_Array_0_block_ram_r_5_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_6_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n955, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n699, q => 
                           load_n_store_RGB_Array_0_block_ram_r_6_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_6_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n956, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n700, q => 
                           load_n_store_RGB_Array_0_block_ram_r_6_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_6_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n957, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n701, q => 
                           load_n_store_RGB_Array_0_block_ram_r_6_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_6_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n958, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n702, q => 
                           load_n_store_RGB_Array_0_block_ram_r_6_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_6_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n959, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n703, q => 
                           load_n_store_RGB_Array_0_block_ram_r_6_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_6_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n960, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n704, q => 
                           load_n_store_RGB_Array_0_block_ram_r_6_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_6_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n961, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n705, q => 
                           load_n_store_RGB_Array_0_block_ram_r_6_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_6_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n962, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n706, q => 
                           load_n_store_RGB_Array_0_block_ram_r_6_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_7_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n963, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n707, q => 
                           load_n_store_RGB_Array_0_block_ram_r_7_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_7_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n964, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n708, q => 
                           load_n_store_RGB_Array_0_block_ram_r_7_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_7_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n965, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n709, q => 
                           load_n_store_RGB_Array_0_block_ram_r_7_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_7_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n966, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n710, q => 
                           load_n_store_RGB_Array_0_block_ram_r_7_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_7_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n967, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n711, q => 
                           load_n_store_RGB_Array_0_block_ram_r_7_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_7_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n968, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n712, q => 
                           load_n_store_RGB_Array_0_block_ram_r_7_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_7_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n969, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n713, q => 
                           load_n_store_RGB_Array_0_block_ram_r_7_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_7_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n970, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n714, q => 
                           load_n_store_RGB_Array_0_block_ram_r_7_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_8_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n971, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n715, q => 
                           load_n_store_RGB_Array_0_block_ram_r_8_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_8_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n972, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n716, q => 
                           load_n_store_RGB_Array_0_block_ram_r_8_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_8_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n973, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n717, q => 
                           load_n_store_RGB_Array_0_block_ram_r_8_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_8_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n974, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n718, q => 
                           load_n_store_RGB_Array_0_block_ram_r_8_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_8_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n975, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n719, q => 
                           load_n_store_RGB_Array_0_block_ram_r_8_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_8_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n976, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n720, q => 
                           load_n_store_RGB_Array_0_block_ram_r_8_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_8_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n977, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n721, q => 
                           load_n_store_RGB_Array_0_block_ram_r_8_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_8_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n978, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n722, q => 
                           load_n_store_RGB_Array_0_block_ram_r_8_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_9_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n979, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n723, q => 
                           load_n_store_RGB_Array_0_block_ram_r_9_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_9_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n980, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n724, q => 
                           load_n_store_RGB_Array_0_block_ram_r_9_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_9_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n981, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n725, q => 
                           load_n_store_RGB_Array_0_block_ram_r_9_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_9_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n982, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n726, q => 
                           load_n_store_RGB_Array_0_block_ram_r_9_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_9_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n983, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n727, q => 
                           load_n_store_RGB_Array_0_block_ram_r_9_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_9_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n984, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n728, q => 
                           load_n_store_RGB_Array_0_block_ram_r_9_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_9_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n985, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n729, q => 
                           load_n_store_RGB_Array_0_block_ram_r_9_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_9_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n986, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n730, q => 
                           load_n_store_RGB_Array_0_block_ram_r_9_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_10_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n987, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n731, q => 
                           load_n_store_RGB_Array_0_block_ram_r_10_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_10_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n988, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n732, q => 
                           load_n_store_RGB_Array_0_block_ram_r_10_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_10_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n989, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n733, q => 
                           load_n_store_RGB_Array_0_block_ram_r_10_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_10_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n990, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n734, q => 
                           load_n_store_RGB_Array_0_block_ram_r_10_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_10_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n991, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n735, q => 
                           load_n_store_RGB_Array_0_block_ram_r_10_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_10_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n992, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n736, q => 
                           load_n_store_RGB_Array_0_block_ram_r_10_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_10_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n993, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n737, q => 
                           load_n_store_RGB_Array_0_block_ram_r_10_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_10_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n994, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n738, q => 
                           load_n_store_RGB_Array_0_block_ram_r_10_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_11_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n995, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n739, q => 
                           load_n_store_RGB_Array_0_block_ram_r_11_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_11_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n996, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n740, q => 
                           load_n_store_RGB_Array_0_block_ram_r_11_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_11_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n997, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n741, q => 
                           load_n_store_RGB_Array_0_block_ram_r_11_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_11_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n998, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n742, q => 
                           load_n_store_RGB_Array_0_block_ram_r_11_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_11_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n999, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n743, q => 
                           load_n_store_RGB_Array_0_block_ram_r_11_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_11_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1000, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n744, q => 
                           load_n_store_RGB_Array_0_block_ram_r_11_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_11_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1001, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n745, q => 
                           load_n_store_RGB_Array_0_block_ram_r_11_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_11_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1002, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n746, q => 
                           load_n_store_RGB_Array_0_block_ram_r_11_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_12_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1003, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n747, q => 
                           load_n_store_RGB_Array_0_block_ram_r_12_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_12_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1004, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n748, q => 
                           load_n_store_RGB_Array_0_block_ram_r_12_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_12_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1005, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n749, q => 
                           load_n_store_RGB_Array_0_block_ram_r_12_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_12_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1006, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n750, q => 
                           load_n_store_RGB_Array_0_block_ram_r_12_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_12_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1007, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n751, q => 
                           load_n_store_RGB_Array_0_block_ram_r_12_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_12_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1008, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n752, q => 
                           load_n_store_RGB_Array_0_block_ram_r_12_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_12_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1009, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n753, q => 
                           load_n_store_RGB_Array_0_block_ram_r_12_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_12_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1010, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n754, q => 
                           load_n_store_RGB_Array_0_block_ram_r_12_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_13_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1011, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n755, q => 
                           load_n_store_RGB_Array_0_block_ram_r_13_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_13_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1012, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n756, q => 
                           load_n_store_RGB_Array_0_block_ram_r_13_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_13_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1013, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n757, q => 
                           load_n_store_RGB_Array_0_block_ram_r_13_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_13_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1014, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n758, q => 
                           load_n_store_RGB_Array_0_block_ram_r_13_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_13_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1015, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n759, q => 
                           load_n_store_RGB_Array_0_block_ram_r_13_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_13_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1016, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n760, q => 
                           load_n_store_RGB_Array_0_block_ram_r_13_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_13_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1017, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n761, q => 
                           load_n_store_RGB_Array_0_block_ram_r_13_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_13_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1018, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n762, q => 
                           load_n_store_RGB_Array_0_block_ram_r_13_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_14_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1019, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n763, q => 
                           load_n_store_RGB_Array_0_block_ram_r_14_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_14_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1020, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n764, q => 
                           load_n_store_RGB_Array_0_block_ram_r_14_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_14_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1021, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n765, q => 
                           load_n_store_RGB_Array_0_block_ram_r_14_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_14_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1022, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n766, q => 
                           load_n_store_RGB_Array_0_block_ram_r_14_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_14_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1023, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n767, q => 
                           load_n_store_RGB_Array_0_block_ram_r_14_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_14_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1024, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n768, q => 
                           load_n_store_RGB_Array_0_block_ram_r_14_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_14_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1025, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n769, q => 
                           load_n_store_RGB_Array_0_block_ram_r_14_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_14_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1026, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n770, q => 
                           load_n_store_RGB_Array_0_block_ram_r_14_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_15_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1027, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n771, q => 
                           load_n_store_RGB_Array_0_block_ram_r_15_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_15_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1028, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n772, q => 
                           load_n_store_RGB_Array_0_block_ram_r_15_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_15_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1029, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n773, q => 
                           load_n_store_RGB_Array_0_block_ram_r_15_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_15_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1030, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n774, q => 
                           load_n_store_RGB_Array_0_block_ram_r_15_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_15_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1031, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n775, q => 
                           load_n_store_RGB_Array_0_block_ram_r_15_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_15_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1032, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n776, q => 
                           load_n_store_RGB_Array_0_block_ram_r_15_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_15_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1033, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n777, q => 
                           load_n_store_RGB_Array_0_block_ram_r_15_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_15_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1034, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n778, q => 
                           load_n_store_RGB_Array_0_block_ram_r_15_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_16_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1035, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n779, q => 
                           load_n_store_RGB_Array_0_block_ram_r_16_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_16_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1036, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n780, q => 
                           load_n_store_RGB_Array_0_block_ram_r_16_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_16_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1037, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n781, q => 
                           load_n_store_RGB_Array_0_block_ram_r_16_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_16_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1038, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n782, q => 
                           load_n_store_RGB_Array_0_block_ram_r_16_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_16_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1039, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n783, q => 
                           load_n_store_RGB_Array_0_block_ram_r_16_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_16_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1040, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n784, q => 
                           load_n_store_RGB_Array_0_block_ram_r_16_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_16_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1041, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n785, q => 
                           load_n_store_RGB_Array_0_block_ram_r_16_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_16_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1042, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n786, q => 
                           load_n_store_RGB_Array_0_block_ram_r_16_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_17_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1043, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n787, q => 
                           load_n_store_RGB_Array_0_block_ram_r_17_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_17_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1044, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n788, q => 
                           load_n_store_RGB_Array_0_block_ram_r_17_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_17_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1045, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n789, q => 
                           load_n_store_RGB_Array_0_block_ram_r_17_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_17_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1046, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n790, q => 
                           load_n_store_RGB_Array_0_block_ram_r_17_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_17_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1047, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n791, q => 
                           load_n_store_RGB_Array_0_block_ram_r_17_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_17_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1048, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n792, q => 
                           load_n_store_RGB_Array_0_block_ram_r_17_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_17_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1049, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n793, q => 
                           load_n_store_RGB_Array_0_block_ram_r_17_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_17_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1050, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n794, q => 
                           load_n_store_RGB_Array_0_block_ram_r_17_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_18_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1051, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n795, q => 
                           load_n_store_RGB_Array_0_block_ram_r_18_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_18_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1052, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n796, q => 
                           load_n_store_RGB_Array_0_block_ram_r_18_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_18_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1053, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n797, q => 
                           load_n_store_RGB_Array_0_block_ram_r_18_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_18_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1054, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n798, q => 
                           load_n_store_RGB_Array_0_block_ram_r_18_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_18_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1055, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n799, q => 
                           load_n_store_RGB_Array_0_block_ram_r_18_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_18_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1056, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n800, q => 
                           load_n_store_RGB_Array_0_block_ram_r_18_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_18_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1057, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n801, q => 
                           load_n_store_RGB_Array_0_block_ram_r_18_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_18_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1058, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n802, q => 
                           load_n_store_RGB_Array_0_block_ram_r_18_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_19_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1059, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n803, q => 
                           load_n_store_RGB_Array_0_block_ram_r_19_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_19_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1060, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n804, q => 
                           load_n_store_RGB_Array_0_block_ram_r_19_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_19_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1061, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n805, q => 
                           load_n_store_RGB_Array_0_block_ram_r_19_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_19_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1062, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n806, q => 
                           load_n_store_RGB_Array_0_block_ram_r_19_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_19_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1063, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n807, q => 
                           load_n_store_RGB_Array_0_block_ram_r_19_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_19_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1064, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n808, q => 
                           load_n_store_RGB_Array_0_block_ram_r_19_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_19_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1065, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n809, q => 
                           load_n_store_RGB_Array_0_block_ram_r_19_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_19_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1066, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n810, q => 
                           load_n_store_RGB_Array_0_block_ram_r_19_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_20_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1067, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n811, q => 
                           load_n_store_RGB_Array_0_block_ram_r_20_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_20_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1068, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n812, q => 
                           load_n_store_RGB_Array_0_block_ram_r_20_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_20_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1069, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n813, q => 
                           load_n_store_RGB_Array_0_block_ram_r_20_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_20_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1070, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n814, q => 
                           load_n_store_RGB_Array_0_block_ram_r_20_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_20_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1071, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n815, q => 
                           load_n_store_RGB_Array_0_block_ram_r_20_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_20_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1072, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n816, q => 
                           load_n_store_RGB_Array_0_block_ram_r_20_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_20_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1073, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n817, q => 
                           load_n_store_RGB_Array_0_block_ram_r_20_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_20_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1074, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n818, q => 
                           load_n_store_RGB_Array_0_block_ram_r_20_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_21_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1075, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n819, q => 
                           load_n_store_RGB_Array_0_block_ram_r_21_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_21_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1076, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n820, q => 
                           load_n_store_RGB_Array_0_block_ram_r_21_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_21_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1077, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n821, q => 
                           load_n_store_RGB_Array_0_block_ram_r_21_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_21_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1078, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n822, q => 
                           load_n_store_RGB_Array_0_block_ram_r_21_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_21_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1079, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n823, q => 
                           load_n_store_RGB_Array_0_block_ram_r_21_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_21_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1080, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n824, q => 
                           load_n_store_RGB_Array_0_block_ram_r_21_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_21_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1081, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n825, q => 
                           load_n_store_RGB_Array_0_block_ram_r_21_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_21_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1082, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n826, q => 
                           load_n_store_RGB_Array_0_block_ram_r_21_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_22_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1083, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n827, q => 
                           load_n_store_RGB_Array_0_block_ram_r_22_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_22_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1084, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n828, q => 
                           load_n_store_RGB_Array_0_block_ram_r_22_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_22_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1085, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n829, q => 
                           load_n_store_RGB_Array_0_block_ram_r_22_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_22_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1086, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n830, q => 
                           load_n_store_RGB_Array_0_block_ram_r_22_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_22_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1087, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n831, q => 
                           load_n_store_RGB_Array_0_block_ram_r_22_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_22_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1088, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n832, q => 
                           load_n_store_RGB_Array_0_block_ram_r_22_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_22_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1089, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n833, q => 
                           load_n_store_RGB_Array_0_block_ram_r_22_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_22_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1090, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n834, q => 
                           load_n_store_RGB_Array_0_block_ram_r_22_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_23_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1091, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n835, q => 
                           load_n_store_RGB_Array_0_block_ram_r_23_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_23_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1092, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n836, q => 
                           load_n_store_RGB_Array_0_block_ram_r_23_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_23_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1093, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n837, q => 
                           load_n_store_RGB_Array_0_block_ram_r_23_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_23_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1094, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n838, q => 
                           load_n_store_RGB_Array_0_block_ram_r_23_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_23_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1095, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n839, q => 
                           load_n_store_RGB_Array_0_block_ram_r_23_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_23_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1096, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n840, q => 
                           load_n_store_RGB_Array_0_block_ram_r_23_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_23_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1097, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n841, q => 
                           load_n_store_RGB_Array_0_block_ram_r_23_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_23_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1098, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n842, q => 
                           load_n_store_RGB_Array_0_block_ram_r_23_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_24_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1099, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n843, q => 
                           load_n_store_RGB_Array_0_block_ram_r_24_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_24_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1100, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n844, q => 
                           load_n_store_RGB_Array_0_block_ram_r_24_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_24_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1101, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n845, q => 
                           load_n_store_RGB_Array_0_block_ram_r_24_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_24_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1102, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n846, q => 
                           load_n_store_RGB_Array_0_block_ram_r_24_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_24_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1103, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n847, q => 
                           load_n_store_RGB_Array_0_block_ram_r_24_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_24_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1104, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n848, q => 
                           load_n_store_RGB_Array_0_block_ram_r_24_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_24_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1105, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n849, q => 
                           load_n_store_RGB_Array_0_block_ram_r_24_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_24_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1106, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n850, q => 
                           load_n_store_RGB_Array_0_block_ram_r_24_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_25_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1107, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n851, q => 
                           load_n_store_RGB_Array_0_block_ram_r_25_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_25_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1108, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n852, q => 
                           load_n_store_RGB_Array_0_block_ram_r_25_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_25_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1109, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n853, q => 
                           load_n_store_RGB_Array_0_block_ram_r_25_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_25_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1110, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n854, q => 
                           load_n_store_RGB_Array_0_block_ram_r_25_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_25_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1111, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n855, q => 
                           load_n_store_RGB_Array_0_block_ram_r_25_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_25_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1112, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n856, q => 
                           load_n_store_RGB_Array_0_block_ram_r_25_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_25_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1113, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n857, q => 
                           load_n_store_RGB_Array_0_block_ram_r_25_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_25_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1114, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n858, q => 
                           load_n_store_RGB_Array_0_block_ram_r_25_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_26_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1115, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n859, q => 
                           load_n_store_RGB_Array_0_block_ram_r_26_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_26_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1116, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n860, q => 
                           load_n_store_RGB_Array_0_block_ram_r_26_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_26_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1117, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n861, q => 
                           load_n_store_RGB_Array_0_block_ram_r_26_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_26_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1118, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n862, q => 
                           load_n_store_RGB_Array_0_block_ram_r_26_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_26_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1119, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n863, q => 
                           load_n_store_RGB_Array_0_block_ram_r_26_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_26_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1120, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n864, q => 
                           load_n_store_RGB_Array_0_block_ram_r_26_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_26_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1121, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n865, q => 
                           load_n_store_RGB_Array_0_block_ram_r_26_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_26_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1122, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n866, q => 
                           load_n_store_RGB_Array_0_block_ram_r_26_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_27_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1123, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n867, q => 
                           load_n_store_RGB_Array_0_block_ram_r_27_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_27_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1124, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n868, q => 
                           load_n_store_RGB_Array_0_block_ram_r_27_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_27_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1125, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n869, q => 
                           load_n_store_RGB_Array_0_block_ram_r_27_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_27_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1126, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n870, q => 
                           load_n_store_RGB_Array_0_block_ram_r_27_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_27_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1127, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n871, q => 
                           load_n_store_RGB_Array_0_block_ram_r_27_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_27_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1128, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n872, q => 
                           load_n_store_RGB_Array_0_block_ram_r_27_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_27_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1129, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n873, q => 
                           load_n_store_RGB_Array_0_block_ram_r_27_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_27_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1130, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n874, q => 
                           load_n_store_RGB_Array_0_block_ram_r_27_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_28_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1131, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n875, q => 
                           load_n_store_RGB_Array_0_block_ram_r_28_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_28_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1132, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n876, q => 
                           load_n_store_RGB_Array_0_block_ram_r_28_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_28_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1133, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n877, q => 
                           load_n_store_RGB_Array_0_block_ram_r_28_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_28_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1134, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n878, q => 
                           load_n_store_RGB_Array_0_block_ram_r_28_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_28_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1135, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n879, q => 
                           load_n_store_RGB_Array_0_block_ram_r_28_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_28_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1136, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n880, q => 
                           load_n_store_RGB_Array_0_block_ram_r_28_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_28_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1137, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n881, q => 
                           load_n_store_RGB_Array_0_block_ram_r_28_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_28_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1138, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n882, q => 
                           load_n_store_RGB_Array_0_block_ram_r_28_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_29_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1139, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n883, q => 
                           load_n_store_RGB_Array_0_block_ram_r_29_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_29_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1140, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n884, q => 
                           load_n_store_RGB_Array_0_block_ram_r_29_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_29_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1141, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n885, q => 
                           load_n_store_RGB_Array_0_block_ram_r_29_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_29_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1142, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n886, q => 
                           load_n_store_RGB_Array_0_block_ram_r_29_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_29_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1143, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n887, q => 
                           load_n_store_RGB_Array_0_block_ram_r_29_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_29_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1144, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n888, q => 
                           load_n_store_RGB_Array_0_block_ram_r_29_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_29_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1145, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n889, q => 
                           load_n_store_RGB_Array_0_block_ram_r_29_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_29_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1146, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n890, q => 
                           load_n_store_RGB_Array_0_block_ram_r_29_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_30_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1147, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n891, q => 
                           load_n_store_RGB_Array_0_block_ram_r_30_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_30_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1148, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n892, q => 
                           load_n_store_RGB_Array_0_block_ram_r_30_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_30_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1149, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n893, q => 
                           load_n_store_RGB_Array_0_block_ram_r_30_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_30_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1150, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n894, q => 
                           load_n_store_RGB_Array_0_block_ram_r_30_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_30_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1151, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n895, q => 
                           load_n_store_RGB_Array_0_block_ram_r_30_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_30_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1152, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n896, q => 
                           load_n_store_RGB_Array_0_block_ram_r_30_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_30_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1153, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n897, q => 
                           load_n_store_RGB_Array_0_block_ram_r_30_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_30_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1154, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n898, q => 
                           load_n_store_RGB_Array_0_block_ram_r_30_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_31_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1155, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n899, q => 
                           load_n_store_RGB_Array_0_block_ram_r_31_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_31_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1156, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n900, q => 
                           load_n_store_RGB_Array_0_block_ram_r_31_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_31_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1157, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n901, q => 
                           load_n_store_RGB_Array_0_block_ram_r_31_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_31_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1158, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n902, q => 
                           load_n_store_RGB_Array_0_block_ram_r_31_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_31_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1159, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n903, q => 
                           load_n_store_RGB_Array_0_block_ram_r_31_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_31_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1160, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n904, q => 
                           load_n_store_RGB_Array_0_block_ram_r_31_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_31_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1161, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n905, q => 
                           load_n_store_RGB_Array_0_block_ram_r_31_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_31_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n1162, gclk => clk, rnot =>
                           load_n_store_RGB_Array_0_n906, q => 
                           load_n_store_RGB_Array_0_block_ram_r_31_7_port);
   n3088 <= '1';
   n3087 <= '1';
   n3086 <= '1';
   n3085 <= '1';
   n3084 <= '1';
   n3083 <= '1';
   n3082 <= '1';
   n3081 <= '1';
   n3080 <= '1';
   n3079 <= '1';
   n3078 <= '1';
   n3077 <= '1';
   n3076 <= '1';
   n3075 <= '1';
   n3074 <= '1';
   n3073 <= '1';
   n3072 <= '1';
   n3071 <= '1';
   n3070 <= '1';
   n3069 <= '1';
   n3068 <= '1';
   n3067 <= '1';
   n3066 <= '1';
   n3065 <= '1';
   n3064 <= '1';
   n3063 <= '1';
   n3062 <= '1';
   n3061 <= '1';
   n3060 <= '1';
   n3059 <= '1';
   n3058 <= '1';
   n3057 <= '1';
   n3056 <= '1';
   n3055 <= '1';
   n3054 <= '1';
   n3053 <= '1';
   n3052 <= '1';
   n3051 <= '1';
   n3050 <= '1';
   n3049 <= '1';
   n3048 <= '1';
   n3047 <= '1';
   n3046 <= '1';
   n3045 <= '1';
   n3044 <= '1';
   n3043 <= '1';
   n3042 <= '1';
   n3041 <= '1';
   n3040 <= '1';
   n3039 <= '1';
   n3038 <= '1';
   n3037 <= '1';
   n3036 <= '1';
   n3035 <= '1';
   n3034 <= '1';
   n3033 <= '1';
   n3032 <= '1';
   n3031 <= '1';
   n3030 <= '1';
   n3029 <= '1';
   n3028 <= '1';
   n3027 <= '1';
   n3026 <= '1';
   n3025 <= '1';
   n3024 <= '1';
   n3023 <= '1';
   n3022 <= '1';
   n3021 <= '1';
   n3020 <= '1';
   n3019 <= '1';
   n3018 <= '1';
   n3017 <= '1';
   n3016 <= '1';
   n3015 <= '1';
   n3014 <= '1';
   n3013 <= '1';
   n3012 <= '1';
   n3011 <= '1';
   n3010 <= '1';
   n3009 <= '1';
   n3008 <= '1';
   n3007 <= '1';
   n3006 <= '1';
   n3005 <= '1';
   n3004 <= '1';
   n3003 <= '1';
   n3002 <= '1';
   n3001 <= '1';
   n3000 <= '1';
   n2999 <= '1';
   n2998 <= '1';
   n2997 <= '1';
   n2996 <= '1';
   n2995 <= '1';
   n2994 <= '1';
   n2993 <= '1';
   n2992 <= '1';
   n2991 <= '1';
   n2990 <= '1';
   n2989 <= '1';
   n2988 <= '1';
   n2987 <= '1';
   n2986 <= '1';
   n2985 <= '1';
   n2984 <= '1';
   n2983 <= '1';
   n2982 <= '1';
   n2981 <= '1';
   n2980 <= '1';
   n2979 <= '1';
   n2978 <= '1';
   n2977 <= '1';
   n2976 <= '1';
   n2975 <= '1';
   n2974 <= '1';
   n2973 <= '1';
   n2972 <= '1';
   n2971 <= '1';
   n2970 <= '1';
   n2969 <= '1';
   n2968 <= '1';
   n2967 <= '1';
   n2966 <= '1';
   n2965 <= '1';
   n2964 <= '1';
   n2963 <= '1';
   n2962 <= '1';
   n2961 <= '1';
   n2960 <= '1';
   n2959 <= '1';
   n2958 <= '1';
   n2957 <= '1';
   n2956 <= '1';
   n2955 <= '1';
   n2954 <= '1';
   n2953 <= '1';
   n2952 <= '1';
   n2951 <= '1';
   n2950 <= '1';
   n2949 <= '1';
   n2948 <= '1';
   n2947 <= '1';
   n2946 <= '1';
   n2945 <= '1';
   n2944 <= '1';
   n2943 <= '1';
   n2942 <= '1';
   n2941 <= '1';
   n2940 <= '1';
   n2939 <= '1';
   n2938 <= '1';
   n2937 <= '1';
   n2936 <= '1';
   n2935 <= '1';
   n2934 <= '1';
   n2933 <= '1';
   n2932 <= '1';
   n2931 <= '1';
   n2930 <= '1';
   n2929 <= '1';
   n2928 <= '1';
   n2927 <= '1';
   n2926 <= '1';
   n2925 <= '1';
   n2924 <= '1';
   n2923 <= '1';
   n2922 <= '1';
   n2921 <= '1';
   n2920 <= '1';
   n2919 <= '1';
   n2918 <= '1';
   n2917 <= '1';
   n2916 <= '1';
   n2915 <= '1';
   n2914 <= '1';
   n2913 <= '1';
   n2912 <= '1';
   n2911 <= '1';
   n2910 <= '1';
   n2909 <= '1';
   n2908 <= '1';
   n2907 <= '1';
   n2906 <= '1';
   n2905 <= '1';
   n2904 <= '1';
   n2903 <= '1';
   n2902 <= '1';
   n2901 <= '1';
   n2900 <= '1';
   n2899 <= '1';
   n2898 <= '1';
   n2897 <= '1';
   n2896 <= '1';
   n2895 <= '1';
   n2894 <= '1';
   n2893 <= '1';
   n2892 <= '1';
   n2891 <= '1';
   n2890 <= '1';
   n2889 <= '1';
   n2888 <= '1';
   n2887 <= '1';
   n2886 <= '1';
   n2885 <= '1';
   n2884 <= '1';
   n2883 <= '1';
   n2882 <= '1';
   n2881 <= '1';
   n2880 <= '1';
   n2879 <= '1';
   n2878 <= '1';
   n2877 <= '1';
   n2876 <= '1';
   n2875 <= '1';
   n2874 <= '1';
   n2873 <= '1';
   n2872 <= '1';
   n2871 <= '1';
   n2870 <= '1';
   n2869 <= '1';
   n2868 <= '1';
   n2867 <= '1';
   n2866 <= '1';
   n2865 <= '1';
   n2864 <= '1';
   n2863 <= '1';
   n2862 <= '1';
   n2861 <= '1';
   n2860 <= '1';
   n2859 <= '1';
   n2858 <= '1';
   n2857 <= '1';
   n2856 <= '1';
   n2855 <= '1';
   n2854 <= '1';
   n2853 <= '1';
   n2852 <= '1';
   n2851 <= '1';
   n2850 <= '1';
   n2849 <= '1';
   n2848 <= '1';
   n2847 <= '1';
   n2846 <= '1';
   n2845 <= '1';
   n2844 <= '1';
   n2843 <= '1';
   n2842 <= '1';
   n2841 <= '1';
   n2840 <= '1';
   n2838 <= '1';
   n2837 <= '1';
   n2835 <= '1';
   n2834 <= '1';
   n2832 <= '1';
   n2831 <= '1';
   n2829 <= '1';
   n2828 <= '1';
   n2826 <= '1';
   n2825 <= '1';
   n2823 <= '1';
   n2822 <= '1';
   n2820 <= '1';
   n2819 <= '1';
   n2817 <= '1';
   load_n_store_RGB_Array_2_data_out_o_reg_0_inst : dff port map( d => n2818, 
                           gclk => clk, rnot => n2817, q => 
                           load_n_store_lazy_out_2_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_0_0_inst : dff port map( d => n3089
                           , gclk => clk, rnot => n2819, q => 
                           load_n_store_RGB_Array_2_block_ram_r_0_0_port);
   load_n_store_RGB_Array_2_data_out_o_reg_1_inst : dff port map( d => n2821, 
                           gclk => clk, rnot => n2820, q => 
                           load_n_store_lazy_out_2_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_0_1_inst : dff port map( d => n3090
                           , gclk => clk, rnot => n2822, q => 
                           load_n_store_RGB_Array_2_block_ram_r_0_1_port);
   load_n_store_RGB_Array_2_data_out_o_reg_2_inst : dff port map( d => n2824, 
                           gclk => clk, rnot => n2823, q => 
                           load_n_store_lazy_out_2_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_0_2_inst : dff port map( d => n3091
                           , gclk => clk, rnot => n2825, q => 
                           load_n_store_RGB_Array_2_block_ram_r_0_2_port);
   load_n_store_RGB_Array_2_data_out_o_reg_3_inst : dff port map( d => n2827, 
                           gclk => clk, rnot => n2826, q => 
                           load_n_store_lazy_out_2_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_0_3_inst : dff port map( d => n3092
                           , gclk => clk, rnot => n2828, q => 
                           load_n_store_RGB_Array_2_block_ram_r_0_3_port);
   load_n_store_RGB_Array_2_data_out_o_reg_4_inst : dff port map( d => n2830, 
                           gclk => clk, rnot => n2829, q => 
                           load_n_store_lazy_out_2_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_0_4_inst : dff port map( d => n3093
                           , gclk => clk, rnot => n2831, q => 
                           load_n_store_RGB_Array_2_block_ram_r_0_4_port);
   load_n_store_RGB_Array_2_data_out_o_reg_5_inst : dff port map( d => n2833, 
                           gclk => clk, rnot => n2832, q => 
                           load_n_store_lazy_out_2_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_0_5_inst : dff port map( d => n3094
                           , gclk => clk, rnot => n2834, q => 
                           load_n_store_RGB_Array_2_block_ram_r_0_5_port);
   load_n_store_RGB_Array_2_data_out_o_reg_6_inst : dff port map( d => n2836, 
                           gclk => clk, rnot => n2835, q => 
                           load_n_store_lazy_out_2_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_0_6_inst : dff port map( d => n3095
                           , gclk => clk, rnot => n2837, q => 
                           load_n_store_RGB_Array_2_block_ram_r_0_6_port);
   load_n_store_RGB_Array_2_data_out_o_reg_7_inst : dff port map( d => n2839, 
                           gclk => clk, rnot => n2838, q => 
                           load_n_store_lazy_out_2_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_0_7_inst : dff port map( d => n3096
                           , gclk => clk, rnot => n2840, q => 
                           load_n_store_RGB_Array_2_block_ram_r_0_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_1_0_inst : dff port map( d => n3097
                           , gclk => clk, rnot => n2841, q => 
                           load_n_store_RGB_Array_2_block_ram_r_1_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_1_1_inst : dff port map( d => n3098
                           , gclk => clk, rnot => n2842, q => 
                           load_n_store_RGB_Array_2_block_ram_r_1_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_1_2_inst : dff port map( d => n3099
                           , gclk => clk, rnot => n2843, q => 
                           load_n_store_RGB_Array_2_block_ram_r_1_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_1_3_inst : dff port map( d => n3100
                           , gclk => clk, rnot => n2844, q => 
                           load_n_store_RGB_Array_2_block_ram_r_1_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_1_4_inst : dff port map( d => n3101
                           , gclk => clk, rnot => n2845, q => 
                           load_n_store_RGB_Array_2_block_ram_r_1_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_1_5_inst : dff port map( d => n3102
                           , gclk => clk, rnot => n2846, q => 
                           load_n_store_RGB_Array_2_block_ram_r_1_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_1_6_inst : dff port map( d => n3103
                           , gclk => clk, rnot => n2847, q => 
                           load_n_store_RGB_Array_2_block_ram_r_1_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_1_7_inst : dff port map( d => n3104
                           , gclk => clk, rnot => n2848, q => 
                           load_n_store_RGB_Array_2_block_ram_r_1_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_2_0_inst : dff port map( d => n3105
                           , gclk => clk, rnot => n2849, q => 
                           load_n_store_RGB_Array_2_block_ram_r_2_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_2_1_inst : dff port map( d => n3106
                           , gclk => clk, rnot => n2850, q => 
                           load_n_store_RGB_Array_2_block_ram_r_2_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_2_2_inst : dff port map( d => n3107
                           , gclk => clk, rnot => n2851, q => 
                           load_n_store_RGB_Array_2_block_ram_r_2_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_2_3_inst : dff port map( d => n3108
                           , gclk => clk, rnot => n2852, q => 
                           load_n_store_RGB_Array_2_block_ram_r_2_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_2_4_inst : dff port map( d => n3109
                           , gclk => clk, rnot => n2853, q => 
                           load_n_store_RGB_Array_2_block_ram_r_2_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_2_5_inst : dff port map( d => n3110
                           , gclk => clk, rnot => n2854, q => 
                           load_n_store_RGB_Array_2_block_ram_r_2_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_2_6_inst : dff port map( d => n3111
                           , gclk => clk, rnot => n2855, q => 
                           load_n_store_RGB_Array_2_block_ram_r_2_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_2_7_inst : dff port map( d => n3112
                           , gclk => clk, rnot => n2856, q => 
                           load_n_store_RGB_Array_2_block_ram_r_2_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_3_0_inst : dff port map( d => n3113
                           , gclk => clk, rnot => n2857, q => 
                           load_n_store_RGB_Array_2_block_ram_r_3_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_3_1_inst : dff port map( d => n3114
                           , gclk => clk, rnot => n2858, q => 
                           load_n_store_RGB_Array_2_block_ram_r_3_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_3_2_inst : dff port map( d => n3115
                           , gclk => clk, rnot => n2859, q => 
                           load_n_store_RGB_Array_2_block_ram_r_3_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_3_3_inst : dff port map( d => n3116
                           , gclk => clk, rnot => n2860, q => 
                           load_n_store_RGB_Array_2_block_ram_r_3_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_3_4_inst : dff port map( d => n3117
                           , gclk => clk, rnot => n2861, q => 
                           load_n_store_RGB_Array_2_block_ram_r_3_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_3_5_inst : dff port map( d => n3118
                           , gclk => clk, rnot => n2862, q => 
                           load_n_store_RGB_Array_2_block_ram_r_3_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_3_6_inst : dff port map( d => n3119
                           , gclk => clk, rnot => n2863, q => 
                           load_n_store_RGB_Array_2_block_ram_r_3_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_3_7_inst : dff port map( d => n3120
                           , gclk => clk, rnot => n2864, q => 
                           load_n_store_RGB_Array_2_block_ram_r_3_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_4_0_inst : dff port map( d => n3121
                           , gclk => clk, rnot => n2865, q => 
                           load_n_store_RGB_Array_2_block_ram_r_4_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_4_1_inst : dff port map( d => n3122
                           , gclk => clk, rnot => n2866, q => 
                           load_n_store_RGB_Array_2_block_ram_r_4_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_4_2_inst : dff port map( d => n3123
                           , gclk => clk, rnot => n2867, q => 
                           load_n_store_RGB_Array_2_block_ram_r_4_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_4_3_inst : dff port map( d => n3124
                           , gclk => clk, rnot => n2868, q => 
                           load_n_store_RGB_Array_2_block_ram_r_4_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_4_4_inst : dff port map( d => n3125
                           , gclk => clk, rnot => n2869, q => 
                           load_n_store_RGB_Array_2_block_ram_r_4_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_4_5_inst : dff port map( d => n3126
                           , gclk => clk, rnot => n2870, q => 
                           load_n_store_RGB_Array_2_block_ram_r_4_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_4_6_inst : dff port map( d => n3127
                           , gclk => clk, rnot => n2871, q => 
                           load_n_store_RGB_Array_2_block_ram_r_4_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_4_7_inst : dff port map( d => n3128
                           , gclk => clk, rnot => n2872, q => 
                           load_n_store_RGB_Array_2_block_ram_r_4_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_5_0_inst : dff port map( d => n3129
                           , gclk => clk, rnot => n2873, q => 
                           load_n_store_RGB_Array_2_block_ram_r_5_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_5_1_inst : dff port map( d => n3130
                           , gclk => clk, rnot => n2874, q => 
                           load_n_store_RGB_Array_2_block_ram_r_5_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_5_2_inst : dff port map( d => n3131
                           , gclk => clk, rnot => n2875, q => 
                           load_n_store_RGB_Array_2_block_ram_r_5_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_5_3_inst : dff port map( d => n3132
                           , gclk => clk, rnot => n2876, q => 
                           load_n_store_RGB_Array_2_block_ram_r_5_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_5_4_inst : dff port map( d => n3133
                           , gclk => clk, rnot => n2877, q => 
                           load_n_store_RGB_Array_2_block_ram_r_5_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_5_5_inst : dff port map( d => n3134
                           , gclk => clk, rnot => n2878, q => 
                           load_n_store_RGB_Array_2_block_ram_r_5_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_5_6_inst : dff port map( d => n3135
                           , gclk => clk, rnot => n2879, q => 
                           load_n_store_RGB_Array_2_block_ram_r_5_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_5_7_inst : dff port map( d => n3136
                           , gclk => clk, rnot => n2880, q => 
                           load_n_store_RGB_Array_2_block_ram_r_5_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_6_0_inst : dff port map( d => n3137
                           , gclk => clk, rnot => n2881, q => 
                           load_n_store_RGB_Array_2_block_ram_r_6_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_6_1_inst : dff port map( d => n3138
                           , gclk => clk, rnot => n2882, q => 
                           load_n_store_RGB_Array_2_block_ram_r_6_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_6_2_inst : dff port map( d => n3139
                           , gclk => clk, rnot => n2883, q => 
                           load_n_store_RGB_Array_2_block_ram_r_6_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_6_3_inst : dff port map( d => n3140
                           , gclk => clk, rnot => n2884, q => 
                           load_n_store_RGB_Array_2_block_ram_r_6_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_6_4_inst : dff port map( d => n3141
                           , gclk => clk, rnot => n2885, q => 
                           load_n_store_RGB_Array_2_block_ram_r_6_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_6_5_inst : dff port map( d => n3142
                           , gclk => clk, rnot => n2886, q => 
                           load_n_store_RGB_Array_2_block_ram_r_6_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_6_6_inst : dff port map( d => n3143
                           , gclk => clk, rnot => n2887, q => 
                           load_n_store_RGB_Array_2_block_ram_r_6_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_6_7_inst : dff port map( d => n3144
                           , gclk => clk, rnot => n2888, q => 
                           load_n_store_RGB_Array_2_block_ram_r_6_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_7_0_inst : dff port map( d => n3145
                           , gclk => clk, rnot => n2889, q => 
                           load_n_store_RGB_Array_2_block_ram_r_7_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_7_1_inst : dff port map( d => n3146
                           , gclk => clk, rnot => n2890, q => 
                           load_n_store_RGB_Array_2_block_ram_r_7_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_7_2_inst : dff port map( d => n3147
                           , gclk => clk, rnot => n2891, q => 
                           load_n_store_RGB_Array_2_block_ram_r_7_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_7_3_inst : dff port map( d => n3148
                           , gclk => clk, rnot => n2892, q => 
                           load_n_store_RGB_Array_2_block_ram_r_7_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_7_4_inst : dff port map( d => n3149
                           , gclk => clk, rnot => n2893, q => 
                           load_n_store_RGB_Array_2_block_ram_r_7_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_7_5_inst : dff port map( d => n3150
                           , gclk => clk, rnot => n2894, q => 
                           load_n_store_RGB_Array_2_block_ram_r_7_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_7_6_inst : dff port map( d => n3151
                           , gclk => clk, rnot => n2895, q => 
                           load_n_store_RGB_Array_2_block_ram_r_7_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_7_7_inst : dff port map( d => n3152
                           , gclk => clk, rnot => n2896, q => 
                           load_n_store_RGB_Array_2_block_ram_r_7_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_8_0_inst : dff port map( d => n3153
                           , gclk => clk, rnot => n2897, q => 
                           load_n_store_RGB_Array_2_block_ram_r_8_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_8_1_inst : dff port map( d => n3154
                           , gclk => clk, rnot => n2898, q => 
                           load_n_store_RGB_Array_2_block_ram_r_8_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_8_2_inst : dff port map( d => n3155
                           , gclk => clk, rnot => n2899, q => 
                           load_n_store_RGB_Array_2_block_ram_r_8_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_8_3_inst : dff port map( d => n3156
                           , gclk => clk, rnot => n2900, q => 
                           load_n_store_RGB_Array_2_block_ram_r_8_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_8_4_inst : dff port map( d => n3157
                           , gclk => clk, rnot => n2901, q => 
                           load_n_store_RGB_Array_2_block_ram_r_8_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_8_5_inst : dff port map( d => n3158
                           , gclk => clk, rnot => n2902, q => 
                           load_n_store_RGB_Array_2_block_ram_r_8_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_8_6_inst : dff port map( d => n3159
                           , gclk => clk, rnot => n2903, q => 
                           load_n_store_RGB_Array_2_block_ram_r_8_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_8_7_inst : dff port map( d => n3160
                           , gclk => clk, rnot => n2904, q => 
                           load_n_store_RGB_Array_2_block_ram_r_8_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_9_0_inst : dff port map( d => n3161
                           , gclk => clk, rnot => n2905, q => 
                           load_n_store_RGB_Array_2_block_ram_r_9_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_9_1_inst : dff port map( d => n3162
                           , gclk => clk, rnot => n2906, q => 
                           load_n_store_RGB_Array_2_block_ram_r_9_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_9_2_inst : dff port map( d => n3163
                           , gclk => clk, rnot => n2907, q => 
                           load_n_store_RGB_Array_2_block_ram_r_9_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_9_3_inst : dff port map( d => n3164
                           , gclk => clk, rnot => n2908, q => 
                           load_n_store_RGB_Array_2_block_ram_r_9_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_9_4_inst : dff port map( d => n3165
                           , gclk => clk, rnot => n2909, q => 
                           load_n_store_RGB_Array_2_block_ram_r_9_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_9_5_inst : dff port map( d => n3166
                           , gclk => clk, rnot => n2910, q => 
                           load_n_store_RGB_Array_2_block_ram_r_9_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_9_6_inst : dff port map( d => n3167
                           , gclk => clk, rnot => n2911, q => 
                           load_n_store_RGB_Array_2_block_ram_r_9_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_9_7_inst : dff port map( d => n3168
                           , gclk => clk, rnot => n2912, q => 
                           load_n_store_RGB_Array_2_block_ram_r_9_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_10_0_inst : dff port map( d => 
                           n3169, gclk => clk, rnot => n2913, q => 
                           load_n_store_RGB_Array_2_block_ram_r_10_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_10_1_inst : dff port map( d => 
                           n3170, gclk => clk, rnot => n2914, q => 
                           load_n_store_RGB_Array_2_block_ram_r_10_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_10_2_inst : dff port map( d => 
                           n3171, gclk => clk, rnot => n2915, q => 
                           load_n_store_RGB_Array_2_block_ram_r_10_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_10_3_inst : dff port map( d => 
                           n3172, gclk => clk, rnot => n2916, q => 
                           load_n_store_RGB_Array_2_block_ram_r_10_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_10_4_inst : dff port map( d => 
                           n3173, gclk => clk, rnot => n2917, q => 
                           load_n_store_RGB_Array_2_block_ram_r_10_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_10_5_inst : dff port map( d => 
                           n3174, gclk => clk, rnot => n2918, q => 
                           load_n_store_RGB_Array_2_block_ram_r_10_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_10_6_inst : dff port map( d => 
                           n3175, gclk => clk, rnot => n2919, q => 
                           load_n_store_RGB_Array_2_block_ram_r_10_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_10_7_inst : dff port map( d => 
                           n3176, gclk => clk, rnot => n2920, q => 
                           load_n_store_RGB_Array_2_block_ram_r_10_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_11_0_inst : dff port map( d => 
                           n3177, gclk => clk, rnot => n2921, q => 
                           load_n_store_RGB_Array_2_block_ram_r_11_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_11_1_inst : dff port map( d => 
                           n3178, gclk => clk, rnot => n2922, q => 
                           load_n_store_RGB_Array_2_block_ram_r_11_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_11_2_inst : dff port map( d => 
                           n3179, gclk => clk, rnot => n2923, q => 
                           load_n_store_RGB_Array_2_block_ram_r_11_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_11_3_inst : dff port map( d => 
                           n3180, gclk => clk, rnot => n2924, q => 
                           load_n_store_RGB_Array_2_block_ram_r_11_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_11_4_inst : dff port map( d => 
                           n3181, gclk => clk, rnot => n2925, q => 
                           load_n_store_RGB_Array_2_block_ram_r_11_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_11_5_inst : dff port map( d => 
                           n3182, gclk => clk, rnot => n2926, q => 
                           load_n_store_RGB_Array_2_block_ram_r_11_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_11_6_inst : dff port map( d => 
                           n3183, gclk => clk, rnot => n2927, q => 
                           load_n_store_RGB_Array_2_block_ram_r_11_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_11_7_inst : dff port map( d => 
                           n3184, gclk => clk, rnot => n2928, q => 
                           load_n_store_RGB_Array_2_block_ram_r_11_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_12_0_inst : dff port map( d => 
                           n3185, gclk => clk, rnot => n2929, q => 
                           load_n_store_RGB_Array_2_block_ram_r_12_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_12_1_inst : dff port map( d => 
                           n3186, gclk => clk, rnot => n2930, q => 
                           load_n_store_RGB_Array_2_block_ram_r_12_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_12_2_inst : dff port map( d => 
                           n3187, gclk => clk, rnot => n2931, q => 
                           load_n_store_RGB_Array_2_block_ram_r_12_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_12_3_inst : dff port map( d => 
                           n3188, gclk => clk, rnot => n2932, q => 
                           load_n_store_RGB_Array_2_block_ram_r_12_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_12_4_inst : dff port map( d => 
                           n3189, gclk => clk, rnot => n2933, q => 
                           load_n_store_RGB_Array_2_block_ram_r_12_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_12_5_inst : dff port map( d => 
                           n3190, gclk => clk, rnot => n2934, q => 
                           load_n_store_RGB_Array_2_block_ram_r_12_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_12_6_inst : dff port map( d => 
                           n3191, gclk => clk, rnot => n2935, q => 
                           load_n_store_RGB_Array_2_block_ram_r_12_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_12_7_inst : dff port map( d => 
                           n3192, gclk => clk, rnot => n2936, q => 
                           load_n_store_RGB_Array_2_block_ram_r_12_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_13_0_inst : dff port map( d => 
                           n3193, gclk => clk, rnot => n2937, q => 
                           load_n_store_RGB_Array_2_block_ram_r_13_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_13_1_inst : dff port map( d => 
                           n3194, gclk => clk, rnot => n2938, q => 
                           load_n_store_RGB_Array_2_block_ram_r_13_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_13_2_inst : dff port map( d => 
                           n3195, gclk => clk, rnot => n2939, q => 
                           load_n_store_RGB_Array_2_block_ram_r_13_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_13_3_inst : dff port map( d => 
                           n3196, gclk => clk, rnot => n2940, q => 
                           load_n_store_RGB_Array_2_block_ram_r_13_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_13_4_inst : dff port map( d => 
                           n3197, gclk => clk, rnot => n2941, q => 
                           load_n_store_RGB_Array_2_block_ram_r_13_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_13_5_inst : dff port map( d => 
                           n3198, gclk => clk, rnot => n2942, q => 
                           load_n_store_RGB_Array_2_block_ram_r_13_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_13_6_inst : dff port map( d => 
                           n3199, gclk => clk, rnot => n2943, q => 
                           load_n_store_RGB_Array_2_block_ram_r_13_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_13_7_inst : dff port map( d => 
                           n3200, gclk => clk, rnot => n2944, q => 
                           load_n_store_RGB_Array_2_block_ram_r_13_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_14_0_inst : dff port map( d => 
                           n3201, gclk => clk, rnot => n2945, q => 
                           load_n_store_RGB_Array_2_block_ram_r_14_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_14_1_inst : dff port map( d => 
                           n3202, gclk => clk, rnot => n2946, q => 
                           load_n_store_RGB_Array_2_block_ram_r_14_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_14_2_inst : dff port map( d => 
                           n3203, gclk => clk, rnot => n2947, q => 
                           load_n_store_RGB_Array_2_block_ram_r_14_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_14_3_inst : dff port map( d => 
                           n3204, gclk => clk, rnot => n2948, q => 
                           load_n_store_RGB_Array_2_block_ram_r_14_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_14_4_inst : dff port map( d => 
                           n3205, gclk => clk, rnot => n2949, q => 
                           load_n_store_RGB_Array_2_block_ram_r_14_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_14_5_inst : dff port map( d => 
                           n3206, gclk => clk, rnot => n2950, q => 
                           load_n_store_RGB_Array_2_block_ram_r_14_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_14_6_inst : dff port map( d => 
                           n3207, gclk => clk, rnot => n2951, q => 
                           load_n_store_RGB_Array_2_block_ram_r_14_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_14_7_inst : dff port map( d => 
                           n3208, gclk => clk, rnot => n2952, q => 
                           load_n_store_RGB_Array_2_block_ram_r_14_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_15_0_inst : dff port map( d => 
                           n3209, gclk => clk, rnot => n2953, q => 
                           load_n_store_RGB_Array_2_block_ram_r_15_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_15_1_inst : dff port map( d => 
                           n3210, gclk => clk, rnot => n2954, q => 
                           load_n_store_RGB_Array_2_block_ram_r_15_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_15_2_inst : dff port map( d => 
                           n3211, gclk => clk, rnot => n2955, q => 
                           load_n_store_RGB_Array_2_block_ram_r_15_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_15_3_inst : dff port map( d => 
                           n3212, gclk => clk, rnot => n2956, q => 
                           load_n_store_RGB_Array_2_block_ram_r_15_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_15_4_inst : dff port map( d => 
                           n3213, gclk => clk, rnot => n2957, q => 
                           load_n_store_RGB_Array_2_block_ram_r_15_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_15_5_inst : dff port map( d => 
                           n3214, gclk => clk, rnot => n2958, q => 
                           load_n_store_RGB_Array_2_block_ram_r_15_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_15_6_inst : dff port map( d => 
                           n3215, gclk => clk, rnot => n2959, q => 
                           load_n_store_RGB_Array_2_block_ram_r_15_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_15_7_inst : dff port map( d => 
                           n3216, gclk => clk, rnot => n2960, q => 
                           load_n_store_RGB_Array_2_block_ram_r_15_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_16_0_inst : dff port map( d => 
                           n3217, gclk => clk, rnot => n2961, q => 
                           load_n_store_RGB_Array_2_block_ram_r_16_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_16_1_inst : dff port map( d => 
                           n3218, gclk => clk, rnot => n2962, q => 
                           load_n_store_RGB_Array_2_block_ram_r_16_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_16_2_inst : dff port map( d => 
                           n3219, gclk => clk, rnot => n2963, q => 
                           load_n_store_RGB_Array_2_block_ram_r_16_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_16_3_inst : dff port map( d => 
                           n3220, gclk => clk, rnot => n2964, q => 
                           load_n_store_RGB_Array_2_block_ram_r_16_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_16_4_inst : dff port map( d => 
                           n3221, gclk => clk, rnot => n2965, q => 
                           load_n_store_RGB_Array_2_block_ram_r_16_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_16_5_inst : dff port map( d => 
                           n3222, gclk => clk, rnot => n2966, q => 
                           load_n_store_RGB_Array_2_block_ram_r_16_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_16_6_inst : dff port map( d => 
                           n3223, gclk => clk, rnot => n2967, q => 
                           load_n_store_RGB_Array_2_block_ram_r_16_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_16_7_inst : dff port map( d => 
                           n3224, gclk => clk, rnot => n2968, q => 
                           load_n_store_RGB_Array_2_block_ram_r_16_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_17_0_inst : dff port map( d => 
                           n3225, gclk => clk, rnot => n2969, q => 
                           load_n_store_RGB_Array_2_block_ram_r_17_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_17_1_inst : dff port map( d => 
                           n3226, gclk => clk, rnot => n2970, q => 
                           load_n_store_RGB_Array_2_block_ram_r_17_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_17_2_inst : dff port map( d => 
                           n3227, gclk => clk, rnot => n2971, q => 
                           load_n_store_RGB_Array_2_block_ram_r_17_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_17_3_inst : dff port map( d => 
                           n3228, gclk => clk, rnot => n2972, q => 
                           load_n_store_RGB_Array_2_block_ram_r_17_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_17_4_inst : dff port map( d => 
                           n3229, gclk => clk, rnot => n2973, q => 
                           load_n_store_RGB_Array_2_block_ram_r_17_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_17_5_inst : dff port map( d => 
                           n3230, gclk => clk, rnot => n2974, q => 
                           load_n_store_RGB_Array_2_block_ram_r_17_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_17_6_inst : dff port map( d => 
                           n3231, gclk => clk, rnot => n2975, q => 
                           load_n_store_RGB_Array_2_block_ram_r_17_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_17_7_inst : dff port map( d => 
                           n3232, gclk => clk, rnot => n2976, q => 
                           load_n_store_RGB_Array_2_block_ram_r_17_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_18_0_inst : dff port map( d => 
                           n3233, gclk => clk, rnot => n2977, q => 
                           load_n_store_RGB_Array_2_block_ram_r_18_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_18_1_inst : dff port map( d => 
                           n3234, gclk => clk, rnot => n2978, q => 
                           load_n_store_RGB_Array_2_block_ram_r_18_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_18_2_inst : dff port map( d => 
                           n3235, gclk => clk, rnot => n2979, q => 
                           load_n_store_RGB_Array_2_block_ram_r_18_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_18_3_inst : dff port map( d => 
                           n3236, gclk => clk, rnot => n2980, q => 
                           load_n_store_RGB_Array_2_block_ram_r_18_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_18_4_inst : dff port map( d => 
                           n3237, gclk => clk, rnot => n2981, q => 
                           load_n_store_RGB_Array_2_block_ram_r_18_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_18_5_inst : dff port map( d => 
                           n3238, gclk => clk, rnot => n2982, q => 
                           load_n_store_RGB_Array_2_block_ram_r_18_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_18_6_inst : dff port map( d => 
                           n3239, gclk => clk, rnot => n2983, q => 
                           load_n_store_RGB_Array_2_block_ram_r_18_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_18_7_inst : dff port map( d => 
                           n3240, gclk => clk, rnot => n2984, q => 
                           load_n_store_RGB_Array_2_block_ram_r_18_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_19_0_inst : dff port map( d => 
                           n3241, gclk => clk, rnot => n2985, q => 
                           load_n_store_RGB_Array_2_block_ram_r_19_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_19_1_inst : dff port map( d => 
                           n3242, gclk => clk, rnot => n2986, q => 
                           load_n_store_RGB_Array_2_block_ram_r_19_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_19_2_inst : dff port map( d => 
                           n3243, gclk => clk, rnot => n2987, q => 
                           load_n_store_RGB_Array_2_block_ram_r_19_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_19_3_inst : dff port map( d => 
                           n3244, gclk => clk, rnot => n2988, q => 
                           load_n_store_RGB_Array_2_block_ram_r_19_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_19_4_inst : dff port map( d => 
                           n3245, gclk => clk, rnot => n2989, q => 
                           load_n_store_RGB_Array_2_block_ram_r_19_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_19_5_inst : dff port map( d => 
                           n3246, gclk => clk, rnot => n2990, q => 
                           load_n_store_RGB_Array_2_block_ram_r_19_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_19_6_inst : dff port map( d => 
                           n3247, gclk => clk, rnot => n2991, q => 
                           load_n_store_RGB_Array_2_block_ram_r_19_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_19_7_inst : dff port map( d => 
                           n3248, gclk => clk, rnot => n2992, q => 
                           load_n_store_RGB_Array_2_block_ram_r_19_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_20_0_inst : dff port map( d => 
                           n3249, gclk => clk, rnot => n2993, q => 
                           load_n_store_RGB_Array_2_block_ram_r_20_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_20_1_inst : dff port map( d => 
                           n3250, gclk => clk, rnot => n2994, q => 
                           load_n_store_RGB_Array_2_block_ram_r_20_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_20_2_inst : dff port map( d => 
                           n3251, gclk => clk, rnot => n2995, q => 
                           load_n_store_RGB_Array_2_block_ram_r_20_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_20_3_inst : dff port map( d => 
                           n3252, gclk => clk, rnot => n2996, q => 
                           load_n_store_RGB_Array_2_block_ram_r_20_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_20_4_inst : dff port map( d => 
                           n3253, gclk => clk, rnot => n2997, q => 
                           load_n_store_RGB_Array_2_block_ram_r_20_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_20_5_inst : dff port map( d => 
                           n3254, gclk => clk, rnot => n2998, q => 
                           load_n_store_RGB_Array_2_block_ram_r_20_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_20_6_inst : dff port map( d => 
                           n3255, gclk => clk, rnot => n2999, q => 
                           load_n_store_RGB_Array_2_block_ram_r_20_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_20_7_inst : dff port map( d => 
                           n3256, gclk => clk, rnot => n3000, q => 
                           load_n_store_RGB_Array_2_block_ram_r_20_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_21_0_inst : dff port map( d => 
                           n3257, gclk => clk, rnot => n3001, q => 
                           load_n_store_RGB_Array_2_block_ram_r_21_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_21_1_inst : dff port map( d => 
                           n3258, gclk => clk, rnot => n3002, q => 
                           load_n_store_RGB_Array_2_block_ram_r_21_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_21_2_inst : dff port map( d => 
                           n3259, gclk => clk, rnot => n3003, q => 
                           load_n_store_RGB_Array_2_block_ram_r_21_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_21_3_inst : dff port map( d => 
                           n3260, gclk => clk, rnot => n3004, q => 
                           load_n_store_RGB_Array_2_block_ram_r_21_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_21_4_inst : dff port map( d => 
                           n3261, gclk => clk, rnot => n3005, q => 
                           load_n_store_RGB_Array_2_block_ram_r_21_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_21_5_inst : dff port map( d => 
                           n3262, gclk => clk, rnot => n3006, q => 
                           load_n_store_RGB_Array_2_block_ram_r_21_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_21_6_inst : dff port map( d => 
                           n3263, gclk => clk, rnot => n3007, q => 
                           load_n_store_RGB_Array_2_block_ram_r_21_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_21_7_inst : dff port map( d => 
                           n3264, gclk => clk, rnot => n3008, q => 
                           load_n_store_RGB_Array_2_block_ram_r_21_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_22_0_inst : dff port map( d => 
                           n3265, gclk => clk, rnot => n3009, q => 
                           load_n_store_RGB_Array_2_block_ram_r_22_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_22_1_inst : dff port map( d => 
                           n3266, gclk => clk, rnot => n3010, q => 
                           load_n_store_RGB_Array_2_block_ram_r_22_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_22_2_inst : dff port map( d => 
                           n3267, gclk => clk, rnot => n3011, q => 
                           load_n_store_RGB_Array_2_block_ram_r_22_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_22_3_inst : dff port map( d => 
                           n3268, gclk => clk, rnot => n3012, q => 
                           load_n_store_RGB_Array_2_block_ram_r_22_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_22_4_inst : dff port map( d => 
                           n3269, gclk => clk, rnot => n3013, q => 
                           load_n_store_RGB_Array_2_block_ram_r_22_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_22_5_inst : dff port map( d => 
                           n3270, gclk => clk, rnot => n3014, q => 
                           load_n_store_RGB_Array_2_block_ram_r_22_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_22_6_inst : dff port map( d => 
                           n3271, gclk => clk, rnot => n3015, q => 
                           load_n_store_RGB_Array_2_block_ram_r_22_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_22_7_inst : dff port map( d => 
                           n3272, gclk => clk, rnot => n3016, q => 
                           load_n_store_RGB_Array_2_block_ram_r_22_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_23_0_inst : dff port map( d => 
                           n3273, gclk => clk, rnot => n3017, q => 
                           load_n_store_RGB_Array_2_block_ram_r_23_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_23_1_inst : dff port map( d => 
                           n3274, gclk => clk, rnot => n3018, q => 
                           load_n_store_RGB_Array_2_block_ram_r_23_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_23_2_inst : dff port map( d => 
                           n3275, gclk => clk, rnot => n3019, q => 
                           load_n_store_RGB_Array_2_block_ram_r_23_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_23_3_inst : dff port map( d => 
                           n3276, gclk => clk, rnot => n3020, q => 
                           load_n_store_RGB_Array_2_block_ram_r_23_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_23_4_inst : dff port map( d => 
                           n3277, gclk => clk, rnot => n3021, q => 
                           load_n_store_RGB_Array_2_block_ram_r_23_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_23_5_inst : dff port map( d => 
                           n3278, gclk => clk, rnot => n3022, q => 
                           load_n_store_RGB_Array_2_block_ram_r_23_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_23_6_inst : dff port map( d => 
                           n3279, gclk => clk, rnot => n3023, q => 
                           load_n_store_RGB_Array_2_block_ram_r_23_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_23_7_inst : dff port map( d => 
                           n3280, gclk => clk, rnot => n3024, q => 
                           load_n_store_RGB_Array_2_block_ram_r_23_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_24_0_inst : dff port map( d => 
                           n3281, gclk => clk, rnot => n3025, q => 
                           load_n_store_RGB_Array_2_block_ram_r_24_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_24_1_inst : dff port map( d => 
                           n3282, gclk => clk, rnot => n3026, q => 
                           load_n_store_RGB_Array_2_block_ram_r_24_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_24_2_inst : dff port map( d => 
                           n3283, gclk => clk, rnot => n3027, q => 
                           load_n_store_RGB_Array_2_block_ram_r_24_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_24_3_inst : dff port map( d => 
                           n3284, gclk => clk, rnot => n3028, q => 
                           load_n_store_RGB_Array_2_block_ram_r_24_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_24_4_inst : dff port map( d => 
                           n3285, gclk => clk, rnot => n3029, q => 
                           load_n_store_RGB_Array_2_block_ram_r_24_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_24_5_inst : dff port map( d => 
                           n3286, gclk => clk, rnot => n3030, q => 
                           load_n_store_RGB_Array_2_block_ram_r_24_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_24_6_inst : dff port map( d => 
                           n3287, gclk => clk, rnot => n3031, q => 
                           load_n_store_RGB_Array_2_block_ram_r_24_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_24_7_inst : dff port map( d => 
                           n3288, gclk => clk, rnot => n3032, q => 
                           load_n_store_RGB_Array_2_block_ram_r_24_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_25_0_inst : dff port map( d => 
                           n3289, gclk => clk, rnot => n3033, q => 
                           load_n_store_RGB_Array_2_block_ram_r_25_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_25_1_inst : dff port map( d => 
                           n3290, gclk => clk, rnot => n3034, q => 
                           load_n_store_RGB_Array_2_block_ram_r_25_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_25_2_inst : dff port map( d => 
                           n3291, gclk => clk, rnot => n3035, q => 
                           load_n_store_RGB_Array_2_block_ram_r_25_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_25_3_inst : dff port map( d => 
                           n3292, gclk => clk, rnot => n3036, q => 
                           load_n_store_RGB_Array_2_block_ram_r_25_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_25_4_inst : dff port map( d => 
                           n3293, gclk => clk, rnot => n3037, q => 
                           load_n_store_RGB_Array_2_block_ram_r_25_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_25_5_inst : dff port map( d => 
                           n3294, gclk => clk, rnot => n3038, q => 
                           load_n_store_RGB_Array_2_block_ram_r_25_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_25_6_inst : dff port map( d => 
                           n3295, gclk => clk, rnot => n3039, q => 
                           load_n_store_RGB_Array_2_block_ram_r_25_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_25_7_inst : dff port map( d => 
                           n3296, gclk => clk, rnot => n3040, q => 
                           load_n_store_RGB_Array_2_block_ram_r_25_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_26_0_inst : dff port map( d => 
                           n3297, gclk => clk, rnot => n3041, q => 
                           load_n_store_RGB_Array_2_block_ram_r_26_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_26_1_inst : dff port map( d => 
                           n3298, gclk => clk, rnot => n3042, q => 
                           load_n_store_RGB_Array_2_block_ram_r_26_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_26_2_inst : dff port map( d => 
                           n3299, gclk => clk, rnot => n3043, q => 
                           load_n_store_RGB_Array_2_block_ram_r_26_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_26_3_inst : dff port map( d => 
                           n3300, gclk => clk, rnot => n3044, q => 
                           load_n_store_RGB_Array_2_block_ram_r_26_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_26_4_inst : dff port map( d => 
                           n3301, gclk => clk, rnot => n3045, q => 
                           load_n_store_RGB_Array_2_block_ram_r_26_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_26_5_inst : dff port map( d => 
                           n3302, gclk => clk, rnot => n3046, q => 
                           load_n_store_RGB_Array_2_block_ram_r_26_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_26_6_inst : dff port map( d => 
                           n3303, gclk => clk, rnot => n3047, q => 
                           load_n_store_RGB_Array_2_block_ram_r_26_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_26_7_inst : dff port map( d => 
                           n3304, gclk => clk, rnot => n3048, q => 
                           load_n_store_RGB_Array_2_block_ram_r_26_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_27_0_inst : dff port map( d => 
                           n3305, gclk => clk, rnot => n3049, q => 
                           load_n_store_RGB_Array_2_block_ram_r_27_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_27_1_inst : dff port map( d => 
                           n3306, gclk => clk, rnot => n3050, q => 
                           load_n_store_RGB_Array_2_block_ram_r_27_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_27_2_inst : dff port map( d => 
                           n3307, gclk => clk, rnot => n3051, q => 
                           load_n_store_RGB_Array_2_block_ram_r_27_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_27_3_inst : dff port map( d => 
                           n3308, gclk => clk, rnot => n3052, q => 
                           load_n_store_RGB_Array_2_block_ram_r_27_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_27_4_inst : dff port map( d => 
                           n3309, gclk => clk, rnot => n3053, q => 
                           load_n_store_RGB_Array_2_block_ram_r_27_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_27_5_inst : dff port map( d => 
                           n3310, gclk => clk, rnot => n3054, q => 
                           load_n_store_RGB_Array_2_block_ram_r_27_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_27_6_inst : dff port map( d => 
                           n3311, gclk => clk, rnot => n3055, q => 
                           load_n_store_RGB_Array_2_block_ram_r_27_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_27_7_inst : dff port map( d => 
                           n3312, gclk => clk, rnot => n3056, q => 
                           load_n_store_RGB_Array_2_block_ram_r_27_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_28_0_inst : dff port map( d => 
                           n3313, gclk => clk, rnot => n3057, q => 
                           load_n_store_RGB_Array_2_block_ram_r_28_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_28_1_inst : dff port map( d => 
                           n3314, gclk => clk, rnot => n3058, q => 
                           load_n_store_RGB_Array_2_block_ram_r_28_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_28_2_inst : dff port map( d => 
                           n3315, gclk => clk, rnot => n3059, q => 
                           load_n_store_RGB_Array_2_block_ram_r_28_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_28_3_inst : dff port map( d => 
                           n3316, gclk => clk, rnot => n3060, q => 
                           load_n_store_RGB_Array_2_block_ram_r_28_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_28_4_inst : dff port map( d => 
                           n3317, gclk => clk, rnot => n3061, q => 
                           load_n_store_RGB_Array_2_block_ram_r_28_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_28_5_inst : dff port map( d => 
                           n3318, gclk => clk, rnot => n3062, q => 
                           load_n_store_RGB_Array_2_block_ram_r_28_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_28_6_inst : dff port map( d => 
                           n3319, gclk => clk, rnot => n3063, q => 
                           load_n_store_RGB_Array_2_block_ram_r_28_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_28_7_inst : dff port map( d => 
                           n3320, gclk => clk, rnot => n3064, q => 
                           load_n_store_RGB_Array_2_block_ram_r_28_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_29_0_inst : dff port map( d => 
                           n3321, gclk => clk, rnot => n3065, q => 
                           load_n_store_RGB_Array_2_block_ram_r_29_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_29_1_inst : dff port map( d => 
                           n3322, gclk => clk, rnot => n3066, q => 
                           load_n_store_RGB_Array_2_block_ram_r_29_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_29_2_inst : dff port map( d => 
                           n3323, gclk => clk, rnot => n3067, q => 
                           load_n_store_RGB_Array_2_block_ram_r_29_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_29_3_inst : dff port map( d => 
                           n3324, gclk => clk, rnot => n3068, q => 
                           load_n_store_RGB_Array_2_block_ram_r_29_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_29_4_inst : dff port map( d => 
                           n3325, gclk => clk, rnot => n3069, q => 
                           load_n_store_RGB_Array_2_block_ram_r_29_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_29_5_inst : dff port map( d => 
                           n3326, gclk => clk, rnot => n3070, q => 
                           load_n_store_RGB_Array_2_block_ram_r_29_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_29_6_inst : dff port map( d => 
                           n3327, gclk => clk, rnot => n3071, q => 
                           load_n_store_RGB_Array_2_block_ram_r_29_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_29_7_inst : dff port map( d => 
                           n3328, gclk => clk, rnot => n3072, q => 
                           load_n_store_RGB_Array_2_block_ram_r_29_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_30_0_inst : dff port map( d => 
                           n3329, gclk => clk, rnot => n3073, q => 
                           load_n_store_RGB_Array_2_block_ram_r_30_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_30_1_inst : dff port map( d => 
                           n3330, gclk => clk, rnot => n3074, q => 
                           load_n_store_RGB_Array_2_block_ram_r_30_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_30_2_inst : dff port map( d => 
                           n3331, gclk => clk, rnot => n3075, q => 
                           load_n_store_RGB_Array_2_block_ram_r_30_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_30_3_inst : dff port map( d => 
                           n3332, gclk => clk, rnot => n3076, q => 
                           load_n_store_RGB_Array_2_block_ram_r_30_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_30_4_inst : dff port map( d => 
                           n3333, gclk => clk, rnot => n3077, q => 
                           load_n_store_RGB_Array_2_block_ram_r_30_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_30_5_inst : dff port map( d => 
                           n3334, gclk => clk, rnot => n3078, q => 
                           load_n_store_RGB_Array_2_block_ram_r_30_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_30_6_inst : dff port map( d => 
                           n3335, gclk => clk, rnot => n3079, q => 
                           load_n_store_RGB_Array_2_block_ram_r_30_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_30_7_inst : dff port map( d => 
                           n3336, gclk => clk, rnot => n3080, q => 
                           load_n_store_RGB_Array_2_block_ram_r_30_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_31_0_inst : dff port map( d => 
                           n3337, gclk => clk, rnot => n3081, q => 
                           load_n_store_RGB_Array_2_block_ram_r_31_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_31_1_inst : dff port map( d => 
                           n3338, gclk => clk, rnot => n3082, q => 
                           load_n_store_RGB_Array_2_block_ram_r_31_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_31_2_inst : dff port map( d => 
                           n3339, gclk => clk, rnot => n3083, q => 
                           load_n_store_RGB_Array_2_block_ram_r_31_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_31_3_inst : dff port map( d => 
                           n3340, gclk => clk, rnot => n3084, q => 
                           load_n_store_RGB_Array_2_block_ram_r_31_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_31_4_inst : dff port map( d => 
                           n3341, gclk => clk, rnot => n3085, q => 
                           load_n_store_RGB_Array_2_block_ram_r_31_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_31_5_inst : dff port map( d => 
                           n3342, gclk => clk, rnot => n3086, q => 
                           load_n_store_RGB_Array_2_block_ram_r_31_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_31_6_inst : dff port map( d => 
                           n3343, gclk => clk, rnot => n3087, q => 
                           load_n_store_RGB_Array_2_block_ram_r_31_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_31_7_inst : dff port map( d => 
                           n3344, gclk => clk, rnot => n3088, q => 
                           load_n_store_RGB_Array_2_block_ram_r_31_7_port);
   n2560 <= '1';
   n2559 <= '1';
   n2558 <= '1';
   n2557 <= '1';
   n2556 <= '1';
   n2555 <= '1';
   n2554 <= '1';
   n2553 <= '1';
   n2552 <= '1';
   n2551 <= '1';
   n2550 <= '1';
   n2549 <= '1';
   n2548 <= '1';
   n2547 <= '1';
   n2546 <= '1';
   n2545 <= '1';
   n2544 <= '1';
   n2543 <= '1';
   n2542 <= '1';
   n2541 <= '1';
   n2540 <= '1';
   n2539 <= '1';
   n2538 <= '1';
   n2537 <= '1';
   n2536 <= '1';
   n2535 <= '1';
   n2534 <= '1';
   n2533 <= '1';
   n2532 <= '1';
   n2531 <= '1';
   n2530 <= '1';
   n2529 <= '1';
   n2528 <= '1';
   n2527 <= '1';
   n2526 <= '1';
   n2525 <= '1';
   n2524 <= '1';
   n2523 <= '1';
   n2522 <= '1';
   n2521 <= '1';
   n2520 <= '1';
   n2519 <= '1';
   n2518 <= '1';
   n2517 <= '1';
   n2516 <= '1';
   n2515 <= '1';
   n2514 <= '1';
   n2513 <= '1';
   n2512 <= '1';
   n2511 <= '1';
   n2510 <= '1';
   n2509 <= '1';
   n2508 <= '1';
   n2507 <= '1';
   n2506 <= '1';
   n2505 <= '1';
   n2504 <= '1';
   n2503 <= '1';
   n2502 <= '1';
   n2501 <= '1';
   n2500 <= '1';
   n2499 <= '1';
   n2498 <= '1';
   n2497 <= '1';
   n2496 <= '1';
   n2495 <= '1';
   n2494 <= '1';
   n2493 <= '1';
   n2492 <= '1';
   n2491 <= '1';
   n2490 <= '1';
   n2489 <= '1';
   n2488 <= '1';
   n2487 <= '1';
   n2486 <= '1';
   n2485 <= '1';
   n2484 <= '1';
   n2483 <= '1';
   n2482 <= '1';
   n2481 <= '1';
   n2480 <= '1';
   n2479 <= '1';
   n2478 <= '1';
   n2477 <= '1';
   n2476 <= '1';
   n2475 <= '1';
   n2474 <= '1';
   n2473 <= '1';
   n2472 <= '1';
   n2471 <= '1';
   n2470 <= '1';
   n2469 <= '1';
   n2468 <= '1';
   n2467 <= '1';
   n2466 <= '1';
   n2465 <= '1';
   n2464 <= '1';
   n2463 <= '1';
   n2462 <= '1';
   n2461 <= '1';
   n2460 <= '1';
   n2459 <= '1';
   n2458 <= '1';
   n2457 <= '1';
   n2456 <= '1';
   n2455 <= '1';
   n2454 <= '1';
   n2453 <= '1';
   n2452 <= '1';
   n2451 <= '1';
   n2450 <= '1';
   n2449 <= '1';
   n2448 <= '1';
   n2447 <= '1';
   n2446 <= '1';
   n2445 <= '1';
   n2444 <= '1';
   n2443 <= '1';
   n2442 <= '1';
   n2441 <= '1';
   n2440 <= '1';
   n2439 <= '1';
   n2438 <= '1';
   n2437 <= '1';
   n2436 <= '1';
   n2435 <= '1';
   n2434 <= '1';
   n2433 <= '1';
   n2432 <= '1';
   n2431 <= '1';
   n2430 <= '1';
   n2429 <= '1';
   n2428 <= '1';
   n2427 <= '1';
   n2426 <= '1';
   n2425 <= '1';
   n2424 <= '1';
   n2423 <= '1';
   n2422 <= '1';
   n2421 <= '1';
   n2420 <= '1';
   n2419 <= '1';
   n2418 <= '1';
   n2417 <= '1';
   n2416 <= '1';
   n2415 <= '1';
   n2414 <= '1';
   n2413 <= '1';
   n2412 <= '1';
   n2411 <= '1';
   n2410 <= '1';
   n2409 <= '1';
   n2408 <= '1';
   n2407 <= '1';
   n2406 <= '1';
   n2405 <= '1';
   n2404 <= '1';
   n2403 <= '1';
   n2402 <= '1';
   n2401 <= '1';
   n2400 <= '1';
   n2399 <= '1';
   n2398 <= '1';
   n2397 <= '1';
   n2396 <= '1';
   n2395 <= '1';
   n2394 <= '1';
   n2393 <= '1';
   n2392 <= '1';
   n2391 <= '1';
   n2390 <= '1';
   n2389 <= '1';
   n2388 <= '1';
   n2387 <= '1';
   n2386 <= '1';
   n2385 <= '1';
   n2384 <= '1';
   n2383 <= '1';
   n2382 <= '1';
   n2381 <= '1';
   n2380 <= '1';
   n2379 <= '1';
   n2378 <= '1';
   n2377 <= '1';
   n2376 <= '1';
   n2375 <= '1';
   n2374 <= '1';
   n2373 <= '1';
   n2372 <= '1';
   n2371 <= '1';
   n2370 <= '1';
   n2369 <= '1';
   n2368 <= '1';
   n2367 <= '1';
   n2366 <= '1';
   n2365 <= '1';
   n2364 <= '1';
   n2363 <= '1';
   n2362 <= '1';
   n2361 <= '1';
   n2360 <= '1';
   n2359 <= '1';
   n2358 <= '1';
   n2357 <= '1';
   n2356 <= '1';
   n2355 <= '1';
   n2354 <= '1';
   n2353 <= '1';
   n2352 <= '1';
   n2351 <= '1';
   n2350 <= '1';
   n2349 <= '1';
   n2348 <= '1';
   n2347 <= '1';
   n2346 <= '1';
   n2345 <= '1';
   n2344 <= '1';
   n2343 <= '1';
   n2342 <= '1';
   n2341 <= '1';
   n2340 <= '1';
   n2339 <= '1';
   n2338 <= '1';
   n2337 <= '1';
   n2336 <= '1';
   n2335 <= '1';
   n2334 <= '1';
   n2333 <= '1';
   n2332 <= '1';
   n2331 <= '1';
   n2330 <= '1';
   n2329 <= '1';
   n2328 <= '1';
   n2327 <= '1';
   n2326 <= '1';
   n2325 <= '1';
   n2324 <= '1';
   n2323 <= '1';
   n2322 <= '1';
   n2321 <= '1';
   n2320 <= '1';
   n2319 <= '1';
   n2318 <= '1';
   n2317 <= '1';
   n2316 <= '1';
   n2315 <= '1';
   n2314 <= '1';
   n2313 <= '1';
   n2312 <= '1';
   n2310 <= '1';
   n2309 <= '1';
   n2307 <= '1';
   n2306 <= '1';
   n2304 <= '1';
   n2303 <= '1';
   n2301 <= '1';
   n2300 <= '1';
   n2298 <= '1';
   n2297 <= '1';
   n2295 <= '1';
   n2294 <= '1';
   n2292 <= '1';
   n2291 <= '1';
   n2289 <= '1';
   load_n_store_RGB_Array_1_data_out_o_reg_0_inst : dff port map( d => n2290, 
                           gclk => clk, rnot => n2289, q => 
                           load_n_store_lazy_out_1_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_0_0_inst : dff port map( d => n2561
                           , gclk => clk, rnot => n2291, q => 
                           load_n_store_RGB_Array_1_block_ram_r_0_0_port);
   load_n_store_RGB_Array_1_data_out_o_reg_1_inst : dff port map( d => n2293, 
                           gclk => clk, rnot => n2292, q => 
                           load_n_store_lazy_out_1_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_0_1_inst : dff port map( d => n2562
                           , gclk => clk, rnot => n2294, q => 
                           load_n_store_RGB_Array_1_block_ram_r_0_1_port);
   load_n_store_RGB_Array_1_data_out_o_reg_2_inst : dff port map( d => n2296, 
                           gclk => clk, rnot => n2295, q => 
                           load_n_store_lazy_out_1_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_0_2_inst : dff port map( d => n2563
                           , gclk => clk, rnot => n2297, q => 
                           load_n_store_RGB_Array_1_block_ram_r_0_2_port);
   load_n_store_RGB_Array_1_data_out_o_reg_3_inst : dff port map( d => n2299, 
                           gclk => clk, rnot => n2298, q => 
                           load_n_store_lazy_out_1_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_0_3_inst : dff port map( d => n2564
                           , gclk => clk, rnot => n2300, q => 
                           load_n_store_RGB_Array_1_block_ram_r_0_3_port);
   load_n_store_RGB_Array_1_data_out_o_reg_4_inst : dff port map( d => n2302, 
                           gclk => clk, rnot => n2301, q => 
                           load_n_store_lazy_out_1_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_0_4_inst : dff port map( d => n2565
                           , gclk => clk, rnot => n2303, q => 
                           load_n_store_RGB_Array_1_block_ram_r_0_4_port);
   load_n_store_RGB_Array_1_data_out_o_reg_5_inst : dff port map( d => n2305, 
                           gclk => clk, rnot => n2304, q => 
                           load_n_store_lazy_out_1_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_0_5_inst : dff port map( d => n2566
                           , gclk => clk, rnot => n2306, q => 
                           load_n_store_RGB_Array_1_block_ram_r_0_5_port);
   load_n_store_RGB_Array_1_data_out_o_reg_6_inst : dff port map( d => n2308, 
                           gclk => clk, rnot => n2307, q => 
                           load_n_store_lazy_out_1_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_0_6_inst : dff port map( d => n2567
                           , gclk => clk, rnot => n2309, q => 
                           load_n_store_RGB_Array_1_block_ram_r_0_6_port);
   load_n_store_RGB_Array_1_data_out_o_reg_7_inst : dff port map( d => n2311, 
                           gclk => clk, rnot => n2310, q => 
                           load_n_store_lazy_out_1_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_0_7_inst : dff port map( d => n2568
                           , gclk => clk, rnot => n2312, q => 
                           load_n_store_RGB_Array_1_block_ram_r_0_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_1_0_inst : dff port map( d => n2569
                           , gclk => clk, rnot => n2313, q => 
                           load_n_store_RGB_Array_1_block_ram_r_1_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_1_1_inst : dff port map( d => n2570
                           , gclk => clk, rnot => n2314, q => 
                           load_n_store_RGB_Array_1_block_ram_r_1_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_1_2_inst : dff port map( d => n2571
                           , gclk => clk, rnot => n2315, q => 
                           load_n_store_RGB_Array_1_block_ram_r_1_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_1_3_inst : dff port map( d => n2572
                           , gclk => clk, rnot => n2316, q => 
                           load_n_store_RGB_Array_1_block_ram_r_1_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_1_4_inst : dff port map( d => n2573
                           , gclk => clk, rnot => n2317, q => 
                           load_n_store_RGB_Array_1_block_ram_r_1_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_1_5_inst : dff port map( d => n2574
                           , gclk => clk, rnot => n2318, q => 
                           load_n_store_RGB_Array_1_block_ram_r_1_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_1_6_inst : dff port map( d => n2575
                           , gclk => clk, rnot => n2319, q => 
                           load_n_store_RGB_Array_1_block_ram_r_1_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_1_7_inst : dff port map( d => n2576
                           , gclk => clk, rnot => n2320, q => 
                           load_n_store_RGB_Array_1_block_ram_r_1_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_2_0_inst : dff port map( d => n2577
                           , gclk => clk, rnot => n2321, q => 
                           load_n_store_RGB_Array_1_block_ram_r_2_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_2_1_inst : dff port map( d => n2578
                           , gclk => clk, rnot => n2322, q => 
                           load_n_store_RGB_Array_1_block_ram_r_2_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_2_2_inst : dff port map( d => n2579
                           , gclk => clk, rnot => n2323, q => 
                           load_n_store_RGB_Array_1_block_ram_r_2_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_2_3_inst : dff port map( d => n2580
                           , gclk => clk, rnot => n2324, q => 
                           load_n_store_RGB_Array_1_block_ram_r_2_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_2_4_inst : dff port map( d => n2581
                           , gclk => clk, rnot => n2325, q => 
                           load_n_store_RGB_Array_1_block_ram_r_2_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_2_5_inst : dff port map( d => n2582
                           , gclk => clk, rnot => n2326, q => 
                           load_n_store_RGB_Array_1_block_ram_r_2_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_2_6_inst : dff port map( d => n2583
                           , gclk => clk, rnot => n2327, q => 
                           load_n_store_RGB_Array_1_block_ram_r_2_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_2_7_inst : dff port map( d => n2584
                           , gclk => clk, rnot => n2328, q => 
                           load_n_store_RGB_Array_1_block_ram_r_2_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_3_0_inst : dff port map( d => n2585
                           , gclk => clk, rnot => n2329, q => 
                           load_n_store_RGB_Array_1_block_ram_r_3_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_3_1_inst : dff port map( d => n2586
                           , gclk => clk, rnot => n2330, q => 
                           load_n_store_RGB_Array_1_block_ram_r_3_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_3_2_inst : dff port map( d => n2587
                           , gclk => clk, rnot => n2331, q => 
                           load_n_store_RGB_Array_1_block_ram_r_3_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_3_3_inst : dff port map( d => n2588
                           , gclk => clk, rnot => n2332, q => 
                           load_n_store_RGB_Array_1_block_ram_r_3_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_3_4_inst : dff port map( d => n2589
                           , gclk => clk, rnot => n2333, q => 
                           load_n_store_RGB_Array_1_block_ram_r_3_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_3_5_inst : dff port map( d => n2590
                           , gclk => clk, rnot => n2334, q => 
                           load_n_store_RGB_Array_1_block_ram_r_3_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_3_6_inst : dff port map( d => n2591
                           , gclk => clk, rnot => n2335, q => 
                           load_n_store_RGB_Array_1_block_ram_r_3_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_3_7_inst : dff port map( d => n2592
                           , gclk => clk, rnot => n2336, q => 
                           load_n_store_RGB_Array_1_block_ram_r_3_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_4_0_inst : dff port map( d => n2593
                           , gclk => clk, rnot => n2337, q => 
                           load_n_store_RGB_Array_1_block_ram_r_4_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_4_1_inst : dff port map( d => n2594
                           , gclk => clk, rnot => n2338, q => 
                           load_n_store_RGB_Array_1_block_ram_r_4_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_4_2_inst : dff port map( d => n2595
                           , gclk => clk, rnot => n2339, q => 
                           load_n_store_RGB_Array_1_block_ram_r_4_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_4_3_inst : dff port map( d => n2596
                           , gclk => clk, rnot => n2340, q => 
                           load_n_store_RGB_Array_1_block_ram_r_4_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_4_4_inst : dff port map( d => n2597
                           , gclk => clk, rnot => n2341, q => 
                           load_n_store_RGB_Array_1_block_ram_r_4_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_4_5_inst : dff port map( d => n2598
                           , gclk => clk, rnot => n2342, q => 
                           load_n_store_RGB_Array_1_block_ram_r_4_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_4_6_inst : dff port map( d => n2599
                           , gclk => clk, rnot => n2343, q => 
                           load_n_store_RGB_Array_1_block_ram_r_4_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_4_7_inst : dff port map( d => n2600
                           , gclk => clk, rnot => n2344, q => 
                           load_n_store_RGB_Array_1_block_ram_r_4_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_5_0_inst : dff port map( d => n2601
                           , gclk => clk, rnot => n2345, q => 
                           load_n_store_RGB_Array_1_block_ram_r_5_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_5_1_inst : dff port map( d => n2602
                           , gclk => clk, rnot => n2346, q => 
                           load_n_store_RGB_Array_1_block_ram_r_5_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_5_2_inst : dff port map( d => n2603
                           , gclk => clk, rnot => n2347, q => 
                           load_n_store_RGB_Array_1_block_ram_r_5_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_5_3_inst : dff port map( d => n2604
                           , gclk => clk, rnot => n2348, q => 
                           load_n_store_RGB_Array_1_block_ram_r_5_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_5_4_inst : dff port map( d => n2605
                           , gclk => clk, rnot => n2349, q => 
                           load_n_store_RGB_Array_1_block_ram_r_5_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_5_5_inst : dff port map( d => n2606
                           , gclk => clk, rnot => n2350, q => 
                           load_n_store_RGB_Array_1_block_ram_r_5_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_5_6_inst : dff port map( d => n2607
                           , gclk => clk, rnot => n2351, q => 
                           load_n_store_RGB_Array_1_block_ram_r_5_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_5_7_inst : dff port map( d => n2608
                           , gclk => clk, rnot => n2352, q => 
                           load_n_store_RGB_Array_1_block_ram_r_5_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_6_0_inst : dff port map( d => n2609
                           , gclk => clk, rnot => n2353, q => 
                           load_n_store_RGB_Array_1_block_ram_r_6_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_6_1_inst : dff port map( d => n2610
                           , gclk => clk, rnot => n2354, q => 
                           load_n_store_RGB_Array_1_block_ram_r_6_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_6_2_inst : dff port map( d => n2611
                           , gclk => clk, rnot => n2355, q => 
                           load_n_store_RGB_Array_1_block_ram_r_6_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_6_3_inst : dff port map( d => n2612
                           , gclk => clk, rnot => n2356, q => 
                           load_n_store_RGB_Array_1_block_ram_r_6_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_6_4_inst : dff port map( d => n2613
                           , gclk => clk, rnot => n2357, q => 
                           load_n_store_RGB_Array_1_block_ram_r_6_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_6_5_inst : dff port map( d => n2614
                           , gclk => clk, rnot => n2358, q => 
                           load_n_store_RGB_Array_1_block_ram_r_6_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_6_6_inst : dff port map( d => n2615
                           , gclk => clk, rnot => n2359, q => 
                           load_n_store_RGB_Array_1_block_ram_r_6_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_6_7_inst : dff port map( d => n2616
                           , gclk => clk, rnot => n2360, q => 
                           load_n_store_RGB_Array_1_block_ram_r_6_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_7_0_inst : dff port map( d => n2617
                           , gclk => clk, rnot => n2361, q => 
                           load_n_store_RGB_Array_1_block_ram_r_7_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_7_1_inst : dff port map( d => n2618
                           , gclk => clk, rnot => n2362, q => 
                           load_n_store_RGB_Array_1_block_ram_r_7_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_7_2_inst : dff port map( d => n2619
                           , gclk => clk, rnot => n2363, q => 
                           load_n_store_RGB_Array_1_block_ram_r_7_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_7_3_inst : dff port map( d => n2620
                           , gclk => clk, rnot => n2364, q => 
                           load_n_store_RGB_Array_1_block_ram_r_7_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_7_4_inst : dff port map( d => n2621
                           , gclk => clk, rnot => n2365, q => 
                           load_n_store_RGB_Array_1_block_ram_r_7_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_7_5_inst : dff port map( d => n2622
                           , gclk => clk, rnot => n2366, q => 
                           load_n_store_RGB_Array_1_block_ram_r_7_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_7_6_inst : dff port map( d => n2623
                           , gclk => clk, rnot => n2367, q => 
                           load_n_store_RGB_Array_1_block_ram_r_7_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_7_7_inst : dff port map( d => n2624
                           , gclk => clk, rnot => n2368, q => 
                           load_n_store_RGB_Array_1_block_ram_r_7_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_8_0_inst : dff port map( d => n2625
                           , gclk => clk, rnot => n2369, q => 
                           load_n_store_RGB_Array_1_block_ram_r_8_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_8_1_inst : dff port map( d => n2626
                           , gclk => clk, rnot => n2370, q => 
                           load_n_store_RGB_Array_1_block_ram_r_8_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_8_2_inst : dff port map( d => n2627
                           , gclk => clk, rnot => n2371, q => 
                           load_n_store_RGB_Array_1_block_ram_r_8_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_8_3_inst : dff port map( d => n2628
                           , gclk => clk, rnot => n2372, q => 
                           load_n_store_RGB_Array_1_block_ram_r_8_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_8_4_inst : dff port map( d => n2629
                           , gclk => clk, rnot => n2373, q => 
                           load_n_store_RGB_Array_1_block_ram_r_8_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_8_5_inst : dff port map( d => n2630
                           , gclk => clk, rnot => n2374, q => 
                           load_n_store_RGB_Array_1_block_ram_r_8_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_8_6_inst : dff port map( d => n2631
                           , gclk => clk, rnot => n2375, q => 
                           load_n_store_RGB_Array_1_block_ram_r_8_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_8_7_inst : dff port map( d => n2632
                           , gclk => clk, rnot => n2376, q => 
                           load_n_store_RGB_Array_1_block_ram_r_8_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_9_0_inst : dff port map( d => n2633
                           , gclk => clk, rnot => n2377, q => 
                           load_n_store_RGB_Array_1_block_ram_r_9_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_9_1_inst : dff port map( d => n2634
                           , gclk => clk, rnot => n2378, q => 
                           load_n_store_RGB_Array_1_block_ram_r_9_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_9_2_inst : dff port map( d => n2635
                           , gclk => clk, rnot => n2379, q => 
                           load_n_store_RGB_Array_1_block_ram_r_9_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_9_3_inst : dff port map( d => n2636
                           , gclk => clk, rnot => n2380, q => 
                           load_n_store_RGB_Array_1_block_ram_r_9_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_9_4_inst : dff port map( d => n2637
                           , gclk => clk, rnot => n2381, q => 
                           load_n_store_RGB_Array_1_block_ram_r_9_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_9_5_inst : dff port map( d => n2638
                           , gclk => clk, rnot => n2382, q => 
                           load_n_store_RGB_Array_1_block_ram_r_9_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_9_6_inst : dff port map( d => n2639
                           , gclk => clk, rnot => n2383, q => 
                           load_n_store_RGB_Array_1_block_ram_r_9_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_9_7_inst : dff port map( d => n2640
                           , gclk => clk, rnot => n2384, q => 
                           load_n_store_RGB_Array_1_block_ram_r_9_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_10_0_inst : dff port map( d => 
                           n2641, gclk => clk, rnot => n2385, q => 
                           load_n_store_RGB_Array_1_block_ram_r_10_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_10_1_inst : dff port map( d => 
                           n2642, gclk => clk, rnot => n2386, q => 
                           load_n_store_RGB_Array_1_block_ram_r_10_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_10_2_inst : dff port map( d => 
                           n2643, gclk => clk, rnot => n2387, q => 
                           load_n_store_RGB_Array_1_block_ram_r_10_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_10_3_inst : dff port map( d => 
                           n2644, gclk => clk, rnot => n2388, q => 
                           load_n_store_RGB_Array_1_block_ram_r_10_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_10_4_inst : dff port map( d => 
                           n2645, gclk => clk, rnot => n2389, q => 
                           load_n_store_RGB_Array_1_block_ram_r_10_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_10_5_inst : dff port map( d => 
                           n2646, gclk => clk, rnot => n2390, q => 
                           load_n_store_RGB_Array_1_block_ram_r_10_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_10_6_inst : dff port map( d => 
                           n2647, gclk => clk, rnot => n2391, q => 
                           load_n_store_RGB_Array_1_block_ram_r_10_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_10_7_inst : dff port map( d => 
                           n2648, gclk => clk, rnot => n2392, q => 
                           load_n_store_RGB_Array_1_block_ram_r_10_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_11_0_inst : dff port map( d => 
                           n2649, gclk => clk, rnot => n2393, q => 
                           load_n_store_RGB_Array_1_block_ram_r_11_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_11_1_inst : dff port map( d => 
                           n2650, gclk => clk, rnot => n2394, q => 
                           load_n_store_RGB_Array_1_block_ram_r_11_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_11_2_inst : dff port map( d => 
                           n2651, gclk => clk, rnot => n2395, q => 
                           load_n_store_RGB_Array_1_block_ram_r_11_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_11_3_inst : dff port map( d => 
                           n2652, gclk => clk, rnot => n2396, q => 
                           load_n_store_RGB_Array_1_block_ram_r_11_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_11_4_inst : dff port map( d => 
                           n2653, gclk => clk, rnot => n2397, q => 
                           load_n_store_RGB_Array_1_block_ram_r_11_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_11_5_inst : dff port map( d => 
                           n2654, gclk => clk, rnot => n2398, q => 
                           load_n_store_RGB_Array_1_block_ram_r_11_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_11_6_inst : dff port map( d => 
                           n2655, gclk => clk, rnot => n2399, q => 
                           load_n_store_RGB_Array_1_block_ram_r_11_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_11_7_inst : dff port map( d => 
                           n2656, gclk => clk, rnot => n2400, q => 
                           load_n_store_RGB_Array_1_block_ram_r_11_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_12_0_inst : dff port map( d => 
                           n2657, gclk => clk, rnot => n2401, q => 
                           load_n_store_RGB_Array_1_block_ram_r_12_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_12_1_inst : dff port map( d => 
                           n2658, gclk => clk, rnot => n2402, q => 
                           load_n_store_RGB_Array_1_block_ram_r_12_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_12_2_inst : dff port map( d => 
                           n2659, gclk => clk, rnot => n2403, q => 
                           load_n_store_RGB_Array_1_block_ram_r_12_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_12_3_inst : dff port map( d => 
                           n2660, gclk => clk, rnot => n2404, q => 
                           load_n_store_RGB_Array_1_block_ram_r_12_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_12_4_inst : dff port map( d => 
                           n2661, gclk => clk, rnot => n2405, q => 
                           load_n_store_RGB_Array_1_block_ram_r_12_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_12_5_inst : dff port map( d => 
                           n2662, gclk => clk, rnot => n2406, q => 
                           load_n_store_RGB_Array_1_block_ram_r_12_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_12_6_inst : dff port map( d => 
                           n2663, gclk => clk, rnot => n2407, q => 
                           load_n_store_RGB_Array_1_block_ram_r_12_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_12_7_inst : dff port map( d => 
                           n2664, gclk => clk, rnot => n2408, q => 
                           load_n_store_RGB_Array_1_block_ram_r_12_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_13_0_inst : dff port map( d => 
                           n2665, gclk => clk, rnot => n2409, q => 
                           load_n_store_RGB_Array_1_block_ram_r_13_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_13_1_inst : dff port map( d => 
                           n2666, gclk => clk, rnot => n2410, q => 
                           load_n_store_RGB_Array_1_block_ram_r_13_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_13_2_inst : dff port map( d => 
                           n2667, gclk => clk, rnot => n2411, q => 
                           load_n_store_RGB_Array_1_block_ram_r_13_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_13_3_inst : dff port map( d => 
                           n2668, gclk => clk, rnot => n2412, q => 
                           load_n_store_RGB_Array_1_block_ram_r_13_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_13_4_inst : dff port map( d => 
                           n2669, gclk => clk, rnot => n2413, q => 
                           load_n_store_RGB_Array_1_block_ram_r_13_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_13_5_inst : dff port map( d => 
                           n2670, gclk => clk, rnot => n2414, q => 
                           load_n_store_RGB_Array_1_block_ram_r_13_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_13_6_inst : dff port map( d => 
                           n2671, gclk => clk, rnot => n2415, q => 
                           load_n_store_RGB_Array_1_block_ram_r_13_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_13_7_inst : dff port map( d => 
                           n2672, gclk => clk, rnot => n2416, q => 
                           load_n_store_RGB_Array_1_block_ram_r_13_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_14_0_inst : dff port map( d => 
                           n2673, gclk => clk, rnot => n2417, q => 
                           load_n_store_RGB_Array_1_block_ram_r_14_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_14_1_inst : dff port map( d => 
                           n2674, gclk => clk, rnot => n2418, q => 
                           load_n_store_RGB_Array_1_block_ram_r_14_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_14_2_inst : dff port map( d => 
                           n2675, gclk => clk, rnot => n2419, q => 
                           load_n_store_RGB_Array_1_block_ram_r_14_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_14_3_inst : dff port map( d => 
                           n2676, gclk => clk, rnot => n2420, q => 
                           load_n_store_RGB_Array_1_block_ram_r_14_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_14_4_inst : dff port map( d => 
                           n2677, gclk => clk, rnot => n2421, q => 
                           load_n_store_RGB_Array_1_block_ram_r_14_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_14_5_inst : dff port map( d => 
                           n2678, gclk => clk, rnot => n2422, q => 
                           load_n_store_RGB_Array_1_block_ram_r_14_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_14_6_inst : dff port map( d => 
                           n2679, gclk => clk, rnot => n2423, q => 
                           load_n_store_RGB_Array_1_block_ram_r_14_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_14_7_inst : dff port map( d => 
                           n2680, gclk => clk, rnot => n2424, q => 
                           load_n_store_RGB_Array_1_block_ram_r_14_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_15_0_inst : dff port map( d => 
                           n2681, gclk => clk, rnot => n2425, q => 
                           load_n_store_RGB_Array_1_block_ram_r_15_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_15_1_inst : dff port map( d => 
                           n2682, gclk => clk, rnot => n2426, q => 
                           load_n_store_RGB_Array_1_block_ram_r_15_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_15_2_inst : dff port map( d => 
                           n2683, gclk => clk, rnot => n2427, q => 
                           load_n_store_RGB_Array_1_block_ram_r_15_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_15_3_inst : dff port map( d => 
                           n2684, gclk => clk, rnot => n2428, q => 
                           load_n_store_RGB_Array_1_block_ram_r_15_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_15_4_inst : dff port map( d => 
                           n2685, gclk => clk, rnot => n2429, q => 
                           load_n_store_RGB_Array_1_block_ram_r_15_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_15_5_inst : dff port map( d => 
                           n2686, gclk => clk, rnot => n2430, q => 
                           load_n_store_RGB_Array_1_block_ram_r_15_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_15_6_inst : dff port map( d => 
                           n2687, gclk => clk, rnot => n2431, q => 
                           load_n_store_RGB_Array_1_block_ram_r_15_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_15_7_inst : dff port map( d => 
                           n2688, gclk => clk, rnot => n2432, q => 
                           load_n_store_RGB_Array_1_block_ram_r_15_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_16_0_inst : dff port map( d => 
                           n2689, gclk => clk, rnot => n2433, q => 
                           load_n_store_RGB_Array_1_block_ram_r_16_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_16_1_inst : dff port map( d => 
                           n2690, gclk => clk, rnot => n2434, q => 
                           load_n_store_RGB_Array_1_block_ram_r_16_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_16_2_inst : dff port map( d => 
                           n2691, gclk => clk, rnot => n2435, q => 
                           load_n_store_RGB_Array_1_block_ram_r_16_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_16_3_inst : dff port map( d => 
                           n2692, gclk => clk, rnot => n2436, q => 
                           load_n_store_RGB_Array_1_block_ram_r_16_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_16_4_inst : dff port map( d => 
                           n2693, gclk => clk, rnot => n2437, q => 
                           load_n_store_RGB_Array_1_block_ram_r_16_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_16_5_inst : dff port map( d => 
                           n2694, gclk => clk, rnot => n2438, q => 
                           load_n_store_RGB_Array_1_block_ram_r_16_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_16_6_inst : dff port map( d => 
                           n2695, gclk => clk, rnot => n2439, q => 
                           load_n_store_RGB_Array_1_block_ram_r_16_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_16_7_inst : dff port map( d => 
                           n2696, gclk => clk, rnot => n2440, q => 
                           load_n_store_RGB_Array_1_block_ram_r_16_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_17_0_inst : dff port map( d => 
                           n2697, gclk => clk, rnot => n2441, q => 
                           load_n_store_RGB_Array_1_block_ram_r_17_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_17_1_inst : dff port map( d => 
                           n2698, gclk => clk, rnot => n2442, q => 
                           load_n_store_RGB_Array_1_block_ram_r_17_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_17_2_inst : dff port map( d => 
                           n2699, gclk => clk, rnot => n2443, q => 
                           load_n_store_RGB_Array_1_block_ram_r_17_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_17_3_inst : dff port map( d => 
                           n2700, gclk => clk, rnot => n2444, q => 
                           load_n_store_RGB_Array_1_block_ram_r_17_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_17_4_inst : dff port map( d => 
                           n2701, gclk => clk, rnot => n2445, q => 
                           load_n_store_RGB_Array_1_block_ram_r_17_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_17_5_inst : dff port map( d => 
                           n2702, gclk => clk, rnot => n2446, q => 
                           load_n_store_RGB_Array_1_block_ram_r_17_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_17_6_inst : dff port map( d => 
                           n2703, gclk => clk, rnot => n2447, q => 
                           load_n_store_RGB_Array_1_block_ram_r_17_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_17_7_inst : dff port map( d => 
                           n2704, gclk => clk, rnot => n2448, q => 
                           load_n_store_RGB_Array_1_block_ram_r_17_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_18_0_inst : dff port map( d => 
                           n2705, gclk => clk, rnot => n2449, q => 
                           load_n_store_RGB_Array_1_block_ram_r_18_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_18_1_inst : dff port map( d => 
                           n2706, gclk => clk, rnot => n2450, q => 
                           load_n_store_RGB_Array_1_block_ram_r_18_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_18_2_inst : dff port map( d => 
                           n2707, gclk => clk, rnot => n2451, q => 
                           load_n_store_RGB_Array_1_block_ram_r_18_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_18_3_inst : dff port map( d => 
                           n2708, gclk => clk, rnot => n2452, q => 
                           load_n_store_RGB_Array_1_block_ram_r_18_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_18_4_inst : dff port map( d => 
                           n2709, gclk => clk, rnot => n2453, q => 
                           load_n_store_RGB_Array_1_block_ram_r_18_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_18_5_inst : dff port map( d => 
                           n2710, gclk => clk, rnot => n2454, q => 
                           load_n_store_RGB_Array_1_block_ram_r_18_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_18_6_inst : dff port map( d => 
                           n2711, gclk => clk, rnot => n2455, q => 
                           load_n_store_RGB_Array_1_block_ram_r_18_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_18_7_inst : dff port map( d => 
                           n2712, gclk => clk, rnot => n2456, q => 
                           load_n_store_RGB_Array_1_block_ram_r_18_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_19_0_inst : dff port map( d => 
                           n2713, gclk => clk, rnot => n2457, q => 
                           load_n_store_RGB_Array_1_block_ram_r_19_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_19_1_inst : dff port map( d => 
                           n2714, gclk => clk, rnot => n2458, q => 
                           load_n_store_RGB_Array_1_block_ram_r_19_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_19_2_inst : dff port map( d => 
                           n2715, gclk => clk, rnot => n2459, q => 
                           load_n_store_RGB_Array_1_block_ram_r_19_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_19_3_inst : dff port map( d => 
                           n2716, gclk => clk, rnot => n2460, q => 
                           load_n_store_RGB_Array_1_block_ram_r_19_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_19_4_inst : dff port map( d => 
                           n2717, gclk => clk, rnot => n2461, q => 
                           load_n_store_RGB_Array_1_block_ram_r_19_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_19_5_inst : dff port map( d => 
                           n2718, gclk => clk, rnot => n2462, q => 
                           load_n_store_RGB_Array_1_block_ram_r_19_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_19_6_inst : dff port map( d => 
                           n2719, gclk => clk, rnot => n2463, q => 
                           load_n_store_RGB_Array_1_block_ram_r_19_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_19_7_inst : dff port map( d => 
                           n2720, gclk => clk, rnot => n2464, q => 
                           load_n_store_RGB_Array_1_block_ram_r_19_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_20_0_inst : dff port map( d => 
                           n2721, gclk => clk, rnot => n2465, q => 
                           load_n_store_RGB_Array_1_block_ram_r_20_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_20_1_inst : dff port map( d => 
                           n2722, gclk => clk, rnot => n2466, q => 
                           load_n_store_RGB_Array_1_block_ram_r_20_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_20_2_inst : dff port map( d => 
                           n2723, gclk => clk, rnot => n2467, q => 
                           load_n_store_RGB_Array_1_block_ram_r_20_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_20_3_inst : dff port map( d => 
                           n2724, gclk => clk, rnot => n2468, q => 
                           load_n_store_RGB_Array_1_block_ram_r_20_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_20_4_inst : dff port map( d => 
                           n2725, gclk => clk, rnot => n2469, q => 
                           load_n_store_RGB_Array_1_block_ram_r_20_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_20_5_inst : dff port map( d => 
                           n2726, gclk => clk, rnot => n2470, q => 
                           load_n_store_RGB_Array_1_block_ram_r_20_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_20_6_inst : dff port map( d => 
                           n2727, gclk => clk, rnot => n2471, q => 
                           load_n_store_RGB_Array_1_block_ram_r_20_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_20_7_inst : dff port map( d => 
                           n2728, gclk => clk, rnot => n2472, q => 
                           load_n_store_RGB_Array_1_block_ram_r_20_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_21_0_inst : dff port map( d => 
                           n2729, gclk => clk, rnot => n2473, q => 
                           load_n_store_RGB_Array_1_block_ram_r_21_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_21_1_inst : dff port map( d => 
                           n2730, gclk => clk, rnot => n2474, q => 
                           load_n_store_RGB_Array_1_block_ram_r_21_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_21_2_inst : dff port map( d => 
                           n2731, gclk => clk, rnot => n2475, q => 
                           load_n_store_RGB_Array_1_block_ram_r_21_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_21_3_inst : dff port map( d => 
                           n2732, gclk => clk, rnot => n2476, q => 
                           load_n_store_RGB_Array_1_block_ram_r_21_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_21_4_inst : dff port map( d => 
                           n2733, gclk => clk, rnot => n2477, q => 
                           load_n_store_RGB_Array_1_block_ram_r_21_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_21_5_inst : dff port map( d => 
                           n2734, gclk => clk, rnot => n2478, q => 
                           load_n_store_RGB_Array_1_block_ram_r_21_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_21_6_inst : dff port map( d => 
                           n2735, gclk => clk, rnot => n2479, q => 
                           load_n_store_RGB_Array_1_block_ram_r_21_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_21_7_inst : dff port map( d => 
                           n2736, gclk => clk, rnot => n2480, q => 
                           load_n_store_RGB_Array_1_block_ram_r_21_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_22_0_inst : dff port map( d => 
                           n2737, gclk => clk, rnot => n2481, q => 
                           load_n_store_RGB_Array_1_block_ram_r_22_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_22_1_inst : dff port map( d => 
                           n2738, gclk => clk, rnot => n2482, q => 
                           load_n_store_RGB_Array_1_block_ram_r_22_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_22_2_inst : dff port map( d => 
                           n2739, gclk => clk, rnot => n2483, q => 
                           load_n_store_RGB_Array_1_block_ram_r_22_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_22_3_inst : dff port map( d => 
                           n2740, gclk => clk, rnot => n2484, q => 
                           load_n_store_RGB_Array_1_block_ram_r_22_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_22_4_inst : dff port map( d => 
                           n2741, gclk => clk, rnot => n2485, q => 
                           load_n_store_RGB_Array_1_block_ram_r_22_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_22_5_inst : dff port map( d => 
                           n2742, gclk => clk, rnot => n2486, q => 
                           load_n_store_RGB_Array_1_block_ram_r_22_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_22_6_inst : dff port map( d => 
                           n2743, gclk => clk, rnot => n2487, q => 
                           load_n_store_RGB_Array_1_block_ram_r_22_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_22_7_inst : dff port map( d => 
                           n2744, gclk => clk, rnot => n2488, q => 
                           load_n_store_RGB_Array_1_block_ram_r_22_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_23_0_inst : dff port map( d => 
                           n2745, gclk => clk, rnot => n2489, q => 
                           load_n_store_RGB_Array_1_block_ram_r_23_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_23_1_inst : dff port map( d => 
                           n2746, gclk => clk, rnot => n2490, q => 
                           load_n_store_RGB_Array_1_block_ram_r_23_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_23_2_inst : dff port map( d => 
                           n2747, gclk => clk, rnot => n2491, q => 
                           load_n_store_RGB_Array_1_block_ram_r_23_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_23_3_inst : dff port map( d => 
                           n2748, gclk => clk, rnot => n2492, q => 
                           load_n_store_RGB_Array_1_block_ram_r_23_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_23_4_inst : dff port map( d => 
                           n2749, gclk => clk, rnot => n2493, q => 
                           load_n_store_RGB_Array_1_block_ram_r_23_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_23_5_inst : dff port map( d => 
                           n2750, gclk => clk, rnot => n2494, q => 
                           load_n_store_RGB_Array_1_block_ram_r_23_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_23_6_inst : dff port map( d => 
                           n2751, gclk => clk, rnot => n2495, q => 
                           load_n_store_RGB_Array_1_block_ram_r_23_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_23_7_inst : dff port map( d => 
                           n2752, gclk => clk, rnot => n2496, q => 
                           load_n_store_RGB_Array_1_block_ram_r_23_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_24_0_inst : dff port map( d => 
                           n2753, gclk => clk, rnot => n2497, q => 
                           load_n_store_RGB_Array_1_block_ram_r_24_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_24_1_inst : dff port map( d => 
                           n2754, gclk => clk, rnot => n2498, q => 
                           load_n_store_RGB_Array_1_block_ram_r_24_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_24_2_inst : dff port map( d => 
                           n2755, gclk => clk, rnot => n2499, q => 
                           load_n_store_RGB_Array_1_block_ram_r_24_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_24_3_inst : dff port map( d => 
                           n2756, gclk => clk, rnot => n2500, q => 
                           load_n_store_RGB_Array_1_block_ram_r_24_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_24_4_inst : dff port map( d => 
                           n2757, gclk => clk, rnot => n2501, q => 
                           load_n_store_RGB_Array_1_block_ram_r_24_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_24_5_inst : dff port map( d => 
                           n2758, gclk => clk, rnot => n2502, q => 
                           load_n_store_RGB_Array_1_block_ram_r_24_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_24_6_inst : dff port map( d => 
                           n2759, gclk => clk, rnot => n2503, q => 
                           load_n_store_RGB_Array_1_block_ram_r_24_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_24_7_inst : dff port map( d => 
                           n2760, gclk => clk, rnot => n2504, q => 
                           load_n_store_RGB_Array_1_block_ram_r_24_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_25_0_inst : dff port map( d => 
                           n2761, gclk => clk, rnot => n2505, q => 
                           load_n_store_RGB_Array_1_block_ram_r_25_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_25_1_inst : dff port map( d => 
                           n2762, gclk => clk, rnot => n2506, q => 
                           load_n_store_RGB_Array_1_block_ram_r_25_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_25_2_inst : dff port map( d => 
                           n2763, gclk => clk, rnot => n2507, q => 
                           load_n_store_RGB_Array_1_block_ram_r_25_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_25_3_inst : dff port map( d => 
                           n2764, gclk => clk, rnot => n2508, q => 
                           load_n_store_RGB_Array_1_block_ram_r_25_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_25_4_inst : dff port map( d => 
                           n2765, gclk => clk, rnot => n2509, q => 
                           load_n_store_RGB_Array_1_block_ram_r_25_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_25_5_inst : dff port map( d => 
                           n2766, gclk => clk, rnot => n2510, q => 
                           load_n_store_RGB_Array_1_block_ram_r_25_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_25_6_inst : dff port map( d => 
                           n2767, gclk => clk, rnot => n2511, q => 
                           load_n_store_RGB_Array_1_block_ram_r_25_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_25_7_inst : dff port map( d => 
                           n2768, gclk => clk, rnot => n2512, q => 
                           load_n_store_RGB_Array_1_block_ram_r_25_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_26_0_inst : dff port map( d => 
                           n2769, gclk => clk, rnot => n2513, q => 
                           load_n_store_RGB_Array_1_block_ram_r_26_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_26_1_inst : dff port map( d => 
                           n2770, gclk => clk, rnot => n2514, q => 
                           load_n_store_RGB_Array_1_block_ram_r_26_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_26_2_inst : dff port map( d => 
                           n2771, gclk => clk, rnot => n2515, q => 
                           load_n_store_RGB_Array_1_block_ram_r_26_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_26_3_inst : dff port map( d => 
                           n2772, gclk => clk, rnot => n2516, q => 
                           load_n_store_RGB_Array_1_block_ram_r_26_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_26_4_inst : dff port map( d => 
                           n2773, gclk => clk, rnot => n2517, q => 
                           load_n_store_RGB_Array_1_block_ram_r_26_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_26_5_inst : dff port map( d => 
                           n2774, gclk => clk, rnot => n2518, q => 
                           load_n_store_RGB_Array_1_block_ram_r_26_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_26_6_inst : dff port map( d => 
                           n2775, gclk => clk, rnot => n2519, q => 
                           load_n_store_RGB_Array_1_block_ram_r_26_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_26_7_inst : dff port map( d => 
                           n2776, gclk => clk, rnot => n2520, q => 
                           load_n_store_RGB_Array_1_block_ram_r_26_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_27_0_inst : dff port map( d => 
                           n2777, gclk => clk, rnot => n2521, q => 
                           load_n_store_RGB_Array_1_block_ram_r_27_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_27_1_inst : dff port map( d => 
                           n2778, gclk => clk, rnot => n2522, q => 
                           load_n_store_RGB_Array_1_block_ram_r_27_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_27_2_inst : dff port map( d => 
                           n2779, gclk => clk, rnot => n2523, q => 
                           load_n_store_RGB_Array_1_block_ram_r_27_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_27_3_inst : dff port map( d => 
                           n2780, gclk => clk, rnot => n2524, q => 
                           load_n_store_RGB_Array_1_block_ram_r_27_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_27_4_inst : dff port map( d => 
                           n2781, gclk => clk, rnot => n2525, q => 
                           load_n_store_RGB_Array_1_block_ram_r_27_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_27_5_inst : dff port map( d => 
                           n2782, gclk => clk, rnot => n2526, q => 
                           load_n_store_RGB_Array_1_block_ram_r_27_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_27_6_inst : dff port map( d => 
                           n2783, gclk => clk, rnot => n2527, q => 
                           load_n_store_RGB_Array_1_block_ram_r_27_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_27_7_inst : dff port map( d => 
                           n2784, gclk => clk, rnot => n2528, q => 
                           load_n_store_RGB_Array_1_block_ram_r_27_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_28_0_inst : dff port map( d => 
                           n2785, gclk => clk, rnot => n2529, q => 
                           load_n_store_RGB_Array_1_block_ram_r_28_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_28_1_inst : dff port map( d => 
                           n2786, gclk => clk, rnot => n2530, q => 
                           load_n_store_RGB_Array_1_block_ram_r_28_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_28_2_inst : dff port map( d => 
                           n2787, gclk => clk, rnot => n2531, q => 
                           load_n_store_RGB_Array_1_block_ram_r_28_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_28_3_inst : dff port map( d => 
                           n2788, gclk => clk, rnot => n2532, q => 
                           load_n_store_RGB_Array_1_block_ram_r_28_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_28_4_inst : dff port map( d => 
                           n2789, gclk => clk, rnot => n2533, q => 
                           load_n_store_RGB_Array_1_block_ram_r_28_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_28_5_inst : dff port map( d => 
                           n2790, gclk => clk, rnot => n2534, q => 
                           load_n_store_RGB_Array_1_block_ram_r_28_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_28_6_inst : dff port map( d => 
                           n2791, gclk => clk, rnot => n2535, q => 
                           load_n_store_RGB_Array_1_block_ram_r_28_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_28_7_inst : dff port map( d => 
                           n2792, gclk => clk, rnot => n2536, q => 
                           load_n_store_RGB_Array_1_block_ram_r_28_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_29_0_inst : dff port map( d => 
                           n2793, gclk => clk, rnot => n2537, q => 
                           load_n_store_RGB_Array_1_block_ram_r_29_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_29_1_inst : dff port map( d => 
                           n2794, gclk => clk, rnot => n2538, q => 
                           load_n_store_RGB_Array_1_block_ram_r_29_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_29_2_inst : dff port map( d => 
                           n2795, gclk => clk, rnot => n2539, q => 
                           load_n_store_RGB_Array_1_block_ram_r_29_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_29_3_inst : dff port map( d => 
                           n2796, gclk => clk, rnot => n2540, q => 
                           load_n_store_RGB_Array_1_block_ram_r_29_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_29_4_inst : dff port map( d => 
                           n2797, gclk => clk, rnot => n2541, q => 
                           load_n_store_RGB_Array_1_block_ram_r_29_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_29_5_inst : dff port map( d => 
                           n2798, gclk => clk, rnot => n2542, q => 
                           load_n_store_RGB_Array_1_block_ram_r_29_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_29_6_inst : dff port map( d => 
                           n2799, gclk => clk, rnot => n2543, q => 
                           load_n_store_RGB_Array_1_block_ram_r_29_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_29_7_inst : dff port map( d => 
                           n2800, gclk => clk, rnot => n2544, q => 
                           load_n_store_RGB_Array_1_block_ram_r_29_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_30_0_inst : dff port map( d => 
                           n2801, gclk => clk, rnot => n2545, q => 
                           load_n_store_RGB_Array_1_block_ram_r_30_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_30_1_inst : dff port map( d => 
                           n2802, gclk => clk, rnot => n2546, q => 
                           load_n_store_RGB_Array_1_block_ram_r_30_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_30_2_inst : dff port map( d => 
                           n2803, gclk => clk, rnot => n2547, q => 
                           load_n_store_RGB_Array_1_block_ram_r_30_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_30_3_inst : dff port map( d => 
                           n2804, gclk => clk, rnot => n2548, q => 
                           load_n_store_RGB_Array_1_block_ram_r_30_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_30_4_inst : dff port map( d => 
                           n2805, gclk => clk, rnot => n2549, q => 
                           load_n_store_RGB_Array_1_block_ram_r_30_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_30_5_inst : dff port map( d => 
                           n2806, gclk => clk, rnot => n2550, q => 
                           load_n_store_RGB_Array_1_block_ram_r_30_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_30_6_inst : dff port map( d => 
                           n2807, gclk => clk, rnot => n2551, q => 
                           load_n_store_RGB_Array_1_block_ram_r_30_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_30_7_inst : dff port map( d => 
                           n2808, gclk => clk, rnot => n2552, q => 
                           load_n_store_RGB_Array_1_block_ram_r_30_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_31_0_inst : dff port map( d => 
                           n2809, gclk => clk, rnot => n2553, q => 
                           load_n_store_RGB_Array_1_block_ram_r_31_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_31_1_inst : dff port map( d => 
                           n2810, gclk => clk, rnot => n2554, q => 
                           load_n_store_RGB_Array_1_block_ram_r_31_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_31_2_inst : dff port map( d => 
                           n2811, gclk => clk, rnot => n2555, q => 
                           load_n_store_RGB_Array_1_block_ram_r_31_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_31_3_inst : dff port map( d => 
                           n2812, gclk => clk, rnot => n2556, q => 
                           load_n_store_RGB_Array_1_block_ram_r_31_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_31_4_inst : dff port map( d => 
                           n2813, gclk => clk, rnot => n2557, q => 
                           load_n_store_RGB_Array_1_block_ram_r_31_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_31_5_inst : dff port map( d => 
                           n2814, gclk => clk, rnot => n2558, q => 
                           load_n_store_RGB_Array_1_block_ram_r_31_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_31_6_inst : dff port map( d => 
                           n2815, gclk => clk, rnot => n2559, q => 
                           load_n_store_RGB_Array_1_block_ram_r_31_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_31_7_inst : dff port map( d => 
                           n2816, gclk => clk, rnot => n2560, q => 
                           load_n_store_RGB_Array_1_block_ram_r_31_7_port);
   U1 : oai22 port map( a => n1, b => n2, c => n3, d => n4, outb => 
                           registers_n296);
   U2 : inv port map( inb => n1, outb => n4);
   U3 : nor2 port map( a => n5, b => n3, outb => n2);
   U4 : oai22 port map( a => n1, b => n6, c => n7, d => n8, outb => 
                           registers_n295);
   U5 : nor2 port map( a => n1, b => registers_s_delay_0_port, outb => n7);
   U6 : aoi12 port map( b => n9, c => n10, a => n11, outb => n1);
   U7 : nand3 port map( a => n12, b => n13, c => n14, outb => registers_n294);
   U8 : inv port map( inb => n11, outb => n12);
   U9 : nand2 port map( a => n15, b => n16, outb => registers_n293);
   U10 : nand3 port map( a => registers_reg_col_inc_1_port, b => 
                           registers_reg_col_inc_0_port, c => n17, outb => n16)
                           ;
   U11 : oai12 port map( b => n18, c => n17, a => registers_reg_col_inc_2_port,
                           outb => n15);
   U12 : inv port map( inb => n19, outb => registers_n292);
   U13 : aoi22 port map( a => addr_i_2_port, b => n20, c => n21, d => 
                           registers_reg_col_inc_2_port, outb => n19);
   U14 : inv port map( inb => n22, outb => registers_n291);
   U15 : aoi22 port map( a => registers_reg_col_inc_0_port, b => n18, c => n23,
                           d => n17, outb => n22);
   U16 : oai22 port map( a => n24, b => n21, c => n20, d => n23, outb => 
                           registers_n290);
   U17 : inv port map( inb => addr_i_0_port, outb => n24);
   U18 : oai12 port map( b => n25, c => n26, a => n27, outb => registers_n289);
   U19 : nand3 port map( a => n17, b => registers_reg_col_inc_0_port, c => n26,
                           outb => n27);
   U20 : aoi12 port map( b => n17, c => n23, a => n18, outb => n25);
   U21 : nor2 port map( a => n28, b => n5, outb => n18);
   U22 : inv port map( inb => registers_reg_col_inc_0_port, outb => n23);
   U23 : oai22 port map( a => n29, b => n21, c => n20, d => n26, outb => 
                           registers_n288);
   U24 : inv port map( inb => registers_reg_col_inc_1_port, outb => n26);
   U25 : inv port map( inb => addr_i_1_port, outb => n29);
   U26 : oai22 port map( a => n30, b => n31, c => n32, d => n33, outb => 
                           registers_n287);
   U27 : nor2 port map( a => n34, b => n35, outb => n32);
   U28 : oai22 port map( a => n36, b => n37, c => registers_reg_cd_0_port, d =>
                           n31, outb => registers_n286);
   U29 : inv port map( inb => n38, outb => registers_n285);
   U30 : aoi12 port map( b => n35, c => n39, a => n40, outb => n38);
   U31 : oai22 port map( a => n41, b => n31, c => n37, d => n42, outb => n40);
   U32 : nand2 port map( a => n35, b => n37, outb => n31);
   U33 : inv port map( inb => n34, outb => n37);
   U34 : nor2 port map( a => n43, b => n11, outb => n34);
   U35 : nor2 port map( a => n44, b => n45, outb => n35);
   U36 : oai12 port map( b => n46, c => n47, a => n48, outb => registers_n284);
   U37 : nand4 port map( a => n5, b => n43, c => registers_reg_row_0_port, d =>
                           n47, outb => n48);
   U38 : aoi12 port map( b => n5, c => n49, a => n50, outb => n46);
   U39 : oai22 port map( a => n51, b => n21, c => n20, d => n47, outb => 
                           registers_n283);
   U40 : inv port map( inb => registers_reg_row_1_port, outb => n47);
   U41 : inv port map( inb => addr_i_4_port, outb => n51);
   U42 : oai12 port map( b => n43, c => n49, a => n52, outb => registers_n282);
   U43 : nand3 port map( a => n5, b => n43, c => n49, outb => n52);
   U44 : inv port map( inb => n50, outb => n43);
   U45 : aoi12 port map( b => n45, c => n11, a => n28, outb => n50);
   U46 : nor2 port map( a => n53, b => n54, outb => n11);
   U47 : oai22 port map( a => n55, b => n21, c => n20, d => n49, outb => 
                           registers_n281);
   U48 : inv port map( inb => registers_reg_row_0_port, outb => n49);
   U49 : inv port map( inb => n20, outb => n21);
   U50 : nor2 port map( a => n28, b => n56, outb => n20);
   U51 : inv port map( inb => addr_i_3_port, outb => n55);
   U52 : nand3 port map( a => n57, b => n58, c => n13, outb => registers_n280);
   U53 : nand3 port map( a => n10, b => n59, c => mem_reg_f, outb => n13);
   U54 : nand2 port map( a => n10, b => n9, outb => n58);
   U55 : nand4 port map( a => n60, b => n44, c => reg_hub_f, d => n61, outb => 
                           n57);
   U56 : oai22 port map( a => n53, b => n62, c => n56, d => n63, outb => 
                           registers_n279);
   U57 : oai12 port map( b => mem_out_b0_7_port, c => n64, a => n65, outb => 
                           n62);
   U58 : aoi22 port map( a => registers_reg_cd_2_port, b => n66, c => n67, d =>
                           n33, outb => n65);
   U59 : inv port map( inb => n68, outb => n67);
   U60 : nor2 port map( a => n69, b => n70, outb => n68);
   U61 : oai22 port map( a => n30, b => mem_out_b0_3_port, c => n71, d => 
                           mem_out_b0_0_port, outb => n70);
   U62 : oai22 port map( a => n72, b => mem_out_b0_2_port, c => n41, d => 
                           mem_out_b0_1_port, outb => n69);
   U63 : oai12 port map( b => mem_out_b0_5_port, c => n41, a => n73, outb => 
                           n66);
   U64 : inv port map( inb => n74, outb => n73);
   U65 : oai22 port map( a => n72, b => mem_out_b0_6_port, c => n71, d => 
                           mem_out_b0_4_port, outb => n74);
   U66 : oai22 port map( a => n61, b => n63, c => n10, d => n75, outb => 
                           registers_n278);
   U67 : inv port map( inb => mem_sipo_b0_7_port, outb => n75);
   U68 : oai22 port map( a => n53, b => n63, c => n56, d => n76, outb => 
                           registers_n277);
   U69 : inv port map( inb => registers_s_mem_sipo_b0_7_port, outb => n63);
   U70 : oai22 port map( a => n61, b => n76, c => n10, d => n77, outb => 
                           registers_n276);
   U71 : inv port map( inb => mem_sipo_b0_6_port, outb => n77);
   U72 : oai22 port map( a => n53, b => n76, c => n56, d => n78, outb => 
                           registers_n275);
   U73 : inv port map( inb => registers_s_mem_sipo_b0_6_port, outb => n76);
   U74 : oai22 port map( a => n61, b => n78, c => n10, d => n79, outb => 
                           registers_n274);
   U75 : inv port map( inb => mem_sipo_b0_5_port, outb => n79);
   U76 : oai22 port map( a => n53, b => n78, c => n56, d => n80, outb => 
                           registers_n273);
   U77 : inv port map( inb => registers_s_mem_sipo_b0_5_port, outb => n78);
   U78 : oai22 port map( a => n61, b => n80, c => n10, d => n81, outb => 
                           registers_n272);
   U79 : inv port map( inb => mem_sipo_b0_4_port, outb => n81);
   U80 : oai22 port map( a => n53, b => n80, c => n56, d => n82, outb => 
                           registers_n271);
   U81 : inv port map( inb => registers_s_mem_sipo_b0_4_port, outb => n80);
   U82 : oai22 port map( a => n61, b => n82, c => n10, d => n83, outb => 
                           registers_n270);
   U83 : inv port map( inb => mem_sipo_b0_3_port, outb => n83);
   U84 : oai22 port map( a => n53, b => n82, c => n56, d => n84, outb => 
                           registers_n269);
   U85 : inv port map( inb => registers_s_mem_sipo_b0_3_port, outb => n82);
   U86 : oai22 port map( a => n61, b => n84, c => n10, d => n85, outb => 
                           registers_n268);
   U87 : inv port map( inb => mem_sipo_b0_2_port, outb => n85);
   U88 : oai22 port map( a => n53, b => n84, c => n56, d => n86, outb => 
                           registers_n267);
   U89 : inv port map( inb => registers_s_mem_sipo_b0_2_port, outb => n84);
   U90 : inv port map( inb => n87, outb => registers_n266);
   U91 : aoi22 port map( a => n10, b => registers_s_mem_sipo_b0_1_port, c => 
                           n61, d => mem_sipo_b0_1_port, outb => n87);
   U92 : oai22 port map( a => n53, b => n86, c => n56, d => n88, outb => 
                           registers_n265);
   U93 : inv port map( inb => registers_s_mem_sipo_b0_1_port, outb => n86);
   U94 : oai22 port map( a => n61, b => n88, c => n10, d => n89, outb => 
                           registers_n264);
   U95 : inv port map( inb => mem_sipo_b0_0_port, outb => n89);
   U96 : inv port map( inb => registers_s_mem_sipo_b0_0_port, outb => n88);
   U97 : oai22 port map( a => n53, b => n90, c => n56, d => n91, outb => 
                           registers_n263);
   U98 : oai12 port map( b => mem_out_r0_7_port, c => n64, a => n92, outb => 
                           n90);
   U99 : aoi22 port map( a => registers_reg_cd_2_port, b => n93, c => n94, d =>
                           n33, outb => n92);
   U100 : inv port map( inb => n95, outb => n94);
   U101 : nor2 port map( a => n96, b => n97, outb => n95);
   U102 : oai22 port map( a => n30, b => mem_out_r0_3_port, c => n71, d => 
                           mem_out_r0_0_port, outb => n97);
   U103 : oai22 port map( a => n72, b => mem_out_r0_2_port, c => n41, d => 
                           mem_out_r0_1_port, outb => n96);
   U104 : oai12 port map( b => mem_out_r0_5_port, c => n41, a => n98, outb => 
                           n93);
   U105 : inv port map( inb => n99, outb => n98);
   U106 : oai22 port map( a => n72, b => mem_out_r0_6_port, c => n71, d => 
                           mem_out_r0_4_port, outb => n99);
   U107 : oai22 port map( a => n53, b => n91, c => n56, d => n100, outb => 
                           registers_n262);
   U108 : oai22 port map( a => n53, b => n100, c => n56, d => n101, outb => 
                           registers_n261);
   U109 : oai22 port map( a => n53, b => n101, c => n56, d => n102, outb => 
                           registers_n260);
   U110 : oai22 port map( a => n53, b => n102, c => n56, d => n103, outb => 
                           registers_n259);
   U111 : oai22 port map( a => n53, b => n103, c => n56, d => n104, outb => 
                           registers_n258);
   U112 : oai22 port map( a => n53, b => n104, c => n56, d => n105, outb => 
                           registers_n257);
   U113 : oai22 port map( a => n53, b => n105, c => n56, d => n106, outb => 
                           registers_n256);
   U114 : inv port map( inb => registers_s_mem_sipo_r0_1_port, outb => n105);
   U115 : oai22 port map( a => n53, b => n107, c => n56, d => n108, outb => 
                           registers_n255);
   U116 : oai12 port map( b => mem_out_g0_7_port, c => n64, a => n109, outb => 
                           n107);
   U117 : aoi22 port map( a => registers_reg_cd_2_port, b => n110, c => n111, d
                           => n33, outb => n109);
   U118 : inv port map( inb => n112, outb => n111);
   U119 : nor2 port map( a => n113, b => n114, outb => n112);
   U120 : oai22 port map( a => n30, b => mem_out_g0_3_port, c => n71, d => 
                           mem_out_g0_0_port, outb => n114);
   U121 : oai22 port map( a => n72, b => mem_out_g0_2_port, c => n41, d => 
                           mem_out_g0_1_port, outb => n113);
   U122 : oai12 port map( b => mem_out_g0_5_port, c => n41, a => n115, outb => 
                           n110);
   U123 : inv port map( inb => n116, outb => n115);
   U124 : oai22 port map( a => n72, b => mem_out_g0_6_port, c => n71, d => 
                           mem_out_g0_4_port, outb => n116);
   U125 : nand2 port map( a => n42, b => n36, outb => n71);
   U126 : inv port map( inb => registers_reg_cd_0_port, outb => n36);
   U127 : inv port map( inb => n39, outb => n72);
   U128 : nor2 port map( a => n42, b => registers_reg_cd_0_port, outb => n39);
   U129 : nand2 port map( a => registers_reg_cd_0_port, b => n42, outb => n41);
   U130 : inv port map( inb => registers_reg_cd_1_port, outb => n42);
   U131 : inv port map( inb => n45, outb => n64);
   U132 : nor2 port map( a => n33, b => n30, outb => n45);
   U133 : nand2 port map( a => registers_reg_cd_1_port, b => 
                           registers_reg_cd_0_port, outb => n30);
   U134 : inv port map( inb => registers_reg_cd_2_port, outb => n33);
   U135 : oai22 port map( a => n53, b => n108, c => n56, d => n117, outb => 
                           registers_n254);
   U136 : oai22 port map( a => n53, b => n117, c => n56, d => n118, outb => 
                           registers_n253);
   U137 : oai22 port map( a => n53, b => n118, c => n56, d => n119, outb => 
                           registers_n252);
   U138 : oai22 port map( a => n53, b => n119, c => n56, d => n120, outb => 
                           registers_n251);
   U139 : oai22 port map( a => n53, b => n120, c => n56, d => n121, outb => 
                           registers_n250);
   U140 : oai22 port map( a => n53, b => n121, c => n56, d => n122, outb => 
                           registers_n249);
   U141 : oai22 port map( a => n53, b => n122, c => n56, d => n123, outb => 
                           registers_n248);
   U142 : inv port map( inb => n53, outb => n56);
   U143 : inv port map( inb => registers_s_mem_sipo_g0_1_port, outb => n122);
   U144 : oai22 port map( a => n61, b => n91, c => n10, d => n124, outb => 
                           registers_n247);
   U145 : inv port map( inb => mem_sipo_r0_7_port, outb => n124);
   U146 : inv port map( inb => registers_s_mem_sipo_r0_7_port, outb => n91);
   U147 : oai22 port map( a => n61, b => n100, c => n10, d => n125, outb => 
                           registers_n246);
   U148 : inv port map( inb => mem_sipo_r0_6_port, outb => n125);
   U149 : inv port map( inb => registers_s_mem_sipo_r0_6_port, outb => n100);
   U150 : oai22 port map( a => n61, b => n101, c => n10, d => n126, outb => 
                           registers_n245);
   U151 : inv port map( inb => mem_sipo_r0_5_port, outb => n126);
   U152 : inv port map( inb => registers_s_mem_sipo_r0_5_port, outb => n101);
   U153 : oai22 port map( a => n61, b => n102, c => n10, d => n127, outb => 
                           registers_n244);
   U154 : inv port map( inb => mem_sipo_r0_4_port, outb => n127);
   U155 : inv port map( inb => registers_s_mem_sipo_r0_4_port, outb => n102);
   U156 : oai22 port map( a => n61, b => n103, c => n10, d => n128, outb => 
                           registers_n243);
   U157 : inv port map( inb => mem_sipo_r0_3_port, outb => n128);
   U158 : inv port map( inb => registers_s_mem_sipo_r0_3_port, outb => n103);
   U159 : oai22 port map( a => n61, b => n104, c => n10, d => n129, outb => 
                           registers_n242);
   U160 : inv port map( inb => mem_sipo_r0_2_port, outb => n129);
   U161 : inv port map( inb => registers_s_mem_sipo_r0_2_port, outb => n104);
   U162 : inv port map( inb => n130, outb => registers_n241);
   U163 : aoi22 port map( a => n10, b => registers_s_mem_sipo_r0_1_port, c => 
                           n61, d => mem_sipo_r0_1_port, outb => n130);
   U164 : oai22 port map( a => n61, b => n106, c => n10, d => n131, outb => 
                           registers_n240);
   U165 : inv port map( inb => mem_sipo_r0_0_port, outb => n131);
   U166 : inv port map( inb => registers_s_mem_sipo_r0_0_port, outb => n106);
   U167 : oai22 port map( a => n61, b => n108, c => n10, d => n132, outb => 
                           registers_n239);
   U168 : inv port map( inb => mem_sipo_g0_7_port, outb => n132);
   U169 : inv port map( inb => registers_s_mem_sipo_g0_7_port, outb => n108);
   U170 : oai22 port map( a => n61, b => n117, c => n10, d => n133, outb => 
                           registers_n238);
   U171 : inv port map( inb => mem_sipo_g0_6_port, outb => n133);
   U172 : inv port map( inb => registers_s_mem_sipo_g0_6_port, outb => n117);
   U173 : oai22 port map( a => n61, b => n118, c => n10, d => n134, outb => 
                           registers_n237);
   U174 : inv port map( inb => mem_sipo_g0_5_port, outb => n134);
   U175 : inv port map( inb => registers_s_mem_sipo_g0_5_port, outb => n118);
   U176 : oai22 port map( a => n61, b => n119, c => n10, d => n135, outb => 
                           registers_n236);
   U177 : inv port map( inb => mem_sipo_g0_4_port, outb => n135);
   U178 : inv port map( inb => registers_s_mem_sipo_g0_4_port, outb => n119);
   U179 : oai22 port map( a => n61, b => n120, c => n10, d => n136, outb => 
                           registers_n235);
   U180 : inv port map( inb => mem_sipo_g0_3_port, outb => n136);
   U181 : inv port map( inb => registers_s_mem_sipo_g0_3_port, outb => n120);
   U182 : oai22 port map( a => n61, b => n121, c => n10, d => n137, outb => 
                           registers_n234);
   U183 : inv port map( inb => mem_sipo_g0_2_port, outb => n137);
   U184 : inv port map( inb => registers_s_mem_sipo_g0_2_port, outb => n121);
   U185 : inv port map( inb => n138, outb => registers_n233);
   U186 : aoi22 port map( a => n10, b => registers_s_mem_sipo_g0_1_port, c => 
                           n61, d => mem_sipo_g0_1_port, outb => n138);
   U187 : oai22 port map( a => n61, b => n123, c => n10, d => n139, outb => 
                           registers_n232);
   U188 : inv port map( inb => mem_sipo_g0_0_port, outb => n139);
   U189 : inv port map( inb => registers_s_mem_sipo_g0_0_port, outb => n123);
   U190 : inv port map( inb => n140, outb => n2218);
   U191 : aoi22 port map( a => n141, b => load_n_store_lazy_out_2_0_port, c => 
                           n142, d => mem_out_r0_0_port, outb => n140);
   U192 : inv port map( inb => n143, outb => n2219);
   U193 : aoi22 port map( a => n141, b => load_n_store_lazy_out_2_1_port, c => 
                           n142, d => mem_out_r0_1_port, outb => n143);
   U194 : inv port map( inb => n144, outb => n2220);
   U195 : aoi22 port map( a => n141, b => load_n_store_lazy_out_2_2_port, c => 
                           n142, d => mem_out_r0_2_port, outb => n144);
   U196 : inv port map( inb => n145, outb => n2221);
   U197 : aoi22 port map( a => n141, b => load_n_store_lazy_out_2_3_port, c => 
                           n142, d => mem_out_r0_3_port, outb => n145);
   U198 : inv port map( inb => n146, outb => n2222);
   U199 : aoi22 port map( a => n141, b => load_n_store_lazy_out_2_4_port, c => 
                           n142, d => mem_out_r0_4_port, outb => n146);
   U200 : inv port map( inb => n147, outb => n2223);
   U201 : aoi22 port map( a => n141, b => load_n_store_lazy_out_2_5_port, c => 
                           n142, d => mem_out_r0_5_port, outb => n147);
   U202 : inv port map( inb => n148, outb => n2224);
   U203 : aoi22 port map( a => n141, b => load_n_store_lazy_out_2_6_port, c => 
                           n142, d => mem_out_r0_6_port, outb => n148);
   U204 : inv port map( inb => n149, outb => n2225);
   U205 : aoi22 port map( a => n141, b => load_n_store_lazy_out_2_7_port, c => 
                           n142, d => mem_out_r0_7_port, outb => n149);
   U206 : inv port map( inb => n150, outb => n2226);
   U207 : aoi22 port map( a => n141, b => load_n_store_lazy_out_1_0_port, c => 
                           n142, d => mem_out_g0_0_port, outb => n150);
   U208 : inv port map( inb => n151, outb => n2227);
   U209 : aoi22 port map( a => n141, b => load_n_store_lazy_out_1_1_port, c => 
                           n142, d => mem_out_g0_1_port, outb => n151);
   U210 : inv port map( inb => n152, outb => n2228);
   U211 : aoi22 port map( a => n141, b => load_n_store_lazy_out_1_2_port, c => 
                           n142, d => mem_out_g0_2_port, outb => n152);
   U212 : inv port map( inb => n153, outb => n2229);
   U213 : aoi22 port map( a => n141, b => load_n_store_lazy_out_1_3_port, c => 
                           n142, d => mem_out_g0_3_port, outb => n153);
   U214 : inv port map( inb => n154, outb => n2230);
   U215 : aoi22 port map( a => n141, b => load_n_store_lazy_out_1_4_port, c => 
                           n142, d => mem_out_g0_4_port, outb => n154);
   U216 : inv port map( inb => n155, outb => n2231);
   U217 : aoi22 port map( a => n141, b => load_n_store_lazy_out_1_5_port, c => 
                           n142, d => mem_out_g0_5_port, outb => n155);
   U218 : inv port map( inb => n156, outb => n2232);
   U219 : aoi22 port map( a => n141, b => load_n_store_lazy_out_1_6_port, c => 
                           n142, d => mem_out_g0_6_port, outb => n156);
   U220 : inv port map( inb => n157, outb => n2233);
   U221 : aoi22 port map( a => n141, b => load_n_store_lazy_out_1_7_port, c => 
                           n142, d => mem_out_g0_7_port, outb => n157);
   U222 : inv port map( inb => n158, outb => n2234);
   U223 : aoi22 port map( a => n141, b => load_n_store_lazy_out_0_0_port, c => 
                           n142, d => mem_out_b0_0_port, outb => n158);
   U224 : inv port map( inb => n159, outb => n2235);
   U225 : aoi22 port map( a => n141, b => load_n_store_lazy_out_0_1_port, c => 
                           n142, d => mem_out_b0_1_port, outb => n159);
   U226 : inv port map( inb => n160, outb => n2236);
   U227 : aoi22 port map( a => n141, b => load_n_store_lazy_out_0_2_port, c => 
                           n142, d => mem_out_b0_2_port, outb => n160);
   U228 : inv port map( inb => n161, outb => n2237);
   U229 : aoi22 port map( a => n141, b => load_n_store_lazy_out_0_3_port, c => 
                           n142, d => mem_out_b0_3_port, outb => n161);
   U230 : inv port map( inb => n162, outb => n2238);
   U231 : aoi22 port map( a => n141, b => load_n_store_lazy_out_0_4_port, c => 
                           n142, d => mem_out_b0_4_port, outb => n162);
   U232 : inv port map( inb => n163, outb => n2239);
   U233 : aoi22 port map( a => n141, b => load_n_store_lazy_out_0_5_port, c => 
                           n142, d => mem_out_b0_5_port, outb => n163);
   U234 : inv port map( inb => n164, outb => n2240);
   U235 : aoi22 port map( a => n141, b => load_n_store_lazy_out_0_6_port, c => 
                           n142, d => mem_out_b0_6_port, outb => n164);
   U236 : inv port map( inb => n165, outb => n2241);
   U237 : aoi22 port map( a => n141, b => load_n_store_lazy_out_0_7_port, c => 
                           n142, d => mem_out_b0_7_port, outb => n165);
   U238 : inv port map( inb => n142, outb => n141);
   U239 : oai22 port map( a => n166, b => n167, c => n168, d => n169, outb => 
                           n2242);
   U240 : inv port map( inb => top_data(16), outb => n167);
   U241 : oai22 port map( a => n166, b => n170, c => n168, d => n171, outb => 
                           n2243);
   U242 : inv port map( inb => top_data(17), outb => n170);
   U243 : oai22 port map( a => n166, b => n172, c => n168, d => n173, outb => 
                           n2244);
   U244 : inv port map( inb => top_data(18), outb => n172);
   U245 : oai22 port map( a => n166, b => n174, c => n168, d => n175, outb => 
                           n2245);
   U246 : inv port map( inb => top_data(19), outb => n174);
   U247 : oai22 port map( a => n166, b => n176, c => n168, d => n177, outb => 
                           n2246);
   U248 : inv port map( inb => top_data(20), outb => n176);
   U249 : oai22 port map( a => n166, b => n178, c => n168, d => n179, outb => 
                           n2247);
   U250 : inv port map( inb => top_data(21), outb => n178);
   U251 : oai22 port map( a => n166, b => n180, c => n168, d => n181, outb => 
                           n2248);
   U252 : inv port map( inb => top_data(22), outb => n180);
   U253 : oai22 port map( a => n166, b => n182, c => n168, d => n183, outb => 
                           n2249);
   U254 : inv port map( inb => top_data(23), outb => n182);
   U255 : oai22 port map( a => n166, b => n184, c => n168, d => n185, outb => 
                           n2250);
   U256 : inv port map( inb => top_data(8), outb => n184);
   U257 : oai22 port map( a => n166, b => n186, c => n168, d => n187, outb => 
                           n2251);
   U258 : inv port map( inb => top_data(9), outb => n186);
   U259 : oai22 port map( a => n166, b => n188, c => n168, d => n189, outb => 
                           n2252);
   U260 : inv port map( inb => top_data(10), outb => n188);
   U261 : oai22 port map( a => n166, b => n190, c => n168, d => n191, outb => 
                           n2253);
   U262 : inv port map( inb => top_data(11), outb => n190);
   U263 : oai22 port map( a => n166, b => n192, c => n168, d => n193, outb => 
                           n2254);
   U264 : inv port map( inb => top_data(12), outb => n192);
   U265 : oai22 port map( a => n166, b => n194, c => n168, d => n195, outb => 
                           n2255);
   U266 : inv port map( inb => top_data(13), outb => n194);
   U267 : oai22 port map( a => n166, b => n196, c => n168, d => n197, outb => 
                           n2256);
   U268 : inv port map( inb => top_data(14), outb => n196);
   U269 : oai22 port map( a => n166, b => n198, c => n168, d => n199, outb => 
                           n2257);
   U270 : inv port map( inb => top_data(15), outb => n198);
   U271 : oai22 port map( a => n166, b => n200, c => n168, d => n201, outb => 
                           n2258);
   U272 : inv port map( inb => top_data(0), outb => n200);
   U273 : oai22 port map( a => n166, b => n202, c => n168, d => n203, outb => 
                           n2259);
   U274 : inv port map( inb => top_data(1), outb => n202);
   U275 : oai22 port map( a => n166, b => n204, c => n168, d => n205, outb => 
                           n2260);
   U276 : inv port map( inb => top_data(2), outb => n204);
   U277 : oai22 port map( a => n166, b => n206, c => n168, d => n207, outb => 
                           n2261);
   U278 : inv port map( inb => top_data(3), outb => n206);
   U279 : oai22 port map( a => n166, b => n208, c => n168, d => n209, outb => 
                           n2262);
   U280 : inv port map( inb => top_data(4), outb => n208);
   U281 : oai22 port map( a => n166, b => n210, c => n168, d => n211, outb => 
                           n2263);
   U282 : inv port map( inb => top_data(5), outb => n210);
   U283 : oai22 port map( a => n166, b => n212, c => n168, d => n213, outb => 
                           n2264);
   U284 : inv port map( inb => top_data(6), outb => n212);
   U285 : oai22 port map( a => n166, b => n214, c => n168, d => n215, outb => 
                           n2265);
   U286 : inv port map( inb => top_data(7), outb => n214);
   U287 : inv port map( inb => n216, outb => n2266);
   U288 : aoi22 port map( a => n217, b => display_out_hub_piso_g0_7_port, c => 
                           n218, d => mem_sipo_g0_7_port, outb => n216);
   U289 : inv port map( inb => n219, outb => n2267);
   U290 : aoi22 port map( a => n217, b => display_out_hub_piso_r0_7_port, c => 
                           n218, d => mem_sipo_r0_7_port, outb => n219);
   U291 : inv port map( inb => n220, outb => n2268);
   U292 : aoi22 port map( a => n217, b => display_out_hub_piso_b0_7_port, c => 
                           n218, d => mem_sipo_b0_7_port, outb => n220);
   U293 : inv port map( inb => n217, outb => n218);
   U294 : inv port map( inb => n221, outb => n2269);
   U295 : aoi22 port map( a => n222, b => n223, c => n224, d => 
                           display_out_clk_timer_6_port, outb => n221);
   U296 : oai12 port map( b => n225, c => n226, a => n227, outb => n224);
   U297 : oai12 port map( b => n227, c => n225, a => n228, outb => n2270);
   U298 : nand4 port map( a => n222, b => n229, c => n230, d => n225, outb => 
                           n228);
   U299 : inv port map( inb => display_out_clk_timer_5_port, outb => n225);
   U300 : aoi12 port map( b => n222, c => display_out_clk_timer_4_port, a => 
                           n231, outb => n227);
   U301 : oai22 port map( a => n226, b => n232, c => n233, d => n234, outb => 
                           n2271);
   U302 : aoi12 port map( b => display_out_clk_timer_0_port, c => n222, a => 
                           n235, outb => n233);
   U303 : oai22 port map( a => n236, b => n237, c => n238, d => n14, outb => 
                           n2272);
   U304 : nor3 port map( a => n239, b => n17, c => n28, outb => n237);
   U305 : nor2 port map( a => n60, b => n240, outb => n28);
   U306 : nor2 port map( a => n53, b => n241, outb => n17);
   U307 : inv port map( inb => n54, outb => n241);
   U308 : nand3 port map( a => registers_reg_col_inc_1_port, b => 
                           registers_reg_col_inc_0_port, c => 
                           registers_reg_col_inc_2_port, outb => n54);
   U309 : nand2 port map( a => mem_reg_f, b => n5, outb => n53);
   U310 : inv port map( inb => n44, outb => n5);
   U311 : nor3 port map( a => n59, b => n61, c => n240, outb => n239);
   U312 : inv port map( inb => n14, outb => n236);
   U313 : nand2 port map( a => n6, b => n60, outb => n14);
   U314 : nand2 port map( a => n242, b => n238, outb => n60);
   U315 : inv port map( inb => registers_mem_to_reg_0_port, outb => n238);
   U316 : inv port map( inb => n243, outb => n6);
   U317 : oai12 port map( b => n61, c => n9, a => n44, outb => n243);
   U318 : nand2 port map( a => registers_mem_to_reg_0_port, b => n242, outb => 
                           n44);
   U319 : nand2 port map( a => n3, b => n8, outb => n9);
   U320 : inv port map( inb => registers_s_delay_1_port, outb => n8);
   U321 : inv port map( inb => registers_s_delay_0_port, outb => n3);
   U322 : inv port map( inb => n10, outb => n61);
   U323 : nor2 port map( a => n242, b => registers_mem_to_reg_0_port, outb => 
                           n10);
   U324 : inv port map( inb => registers_mem_to_reg_1_port, outb => n242);
   U325 : oai22 port map( a => n244, b => n245, c => n246, d => n247, outb => 
                           n2273);
   U326 : aoi12 port map( b => display_out_disp_timer_30_port, c => n248, a => 
                           n249, outb => n246);
   U327 : inv port map( inb => n250, outb => n2274);
   U328 : aoi12 port map( b => n249, c => display_out_disp_timer_30_port, a => 
                           n251, outb => n250);
   U329 : nor3 port map( a => n252, b => display_out_disp_timer_29_port, c => 
                           display_out_disp_timer_30_port, outb => n251);
   U330 : oai12 port map( b => n244, c => n253, a => n254, outb => n249);
   U331 : oai22 port map( a => n254, b => n253, c => 
                           display_out_disp_timer_29_port, d => n252, outb => 
                           n2275);
   U332 : aoi12 port map( b => n248, c => n255, a => n256, outb => n254);
   U333 : oai12 port map( b => n257, c => n258, a => n252, outb => n2276);
   U334 : nand2 port map( a => n259, b => n248, outb => n252);
   U335 : aoi12 port map( b => display_out_disp_timer_27_port, c => n248, a => 
                           n260, outb => n257);
   U336 : oai12 port map( b => n261, c => n262, a => n263, outb => n2277);
   U337 : nand3 port map( a => n264, b => n248, c => n262, outb => n263);
   U338 : inv port map( inb => n260, outb => n261);
   U339 : oai12 port map( b => n244, c => n264, a => n265, outb => n260);
   U340 : inv port map( inb => n266, outb => n2278);
   U341 : aoi22 port map( a => n248, b => n264, c => n267, d => 
                           display_out_disp_timer_26_port, outb => n266);
   U342 : oai12 port map( b => n268, c => n244, a => n269, outb => n267);
   U343 : oai12 port map( b => n269, c => n268, a => n270, outb => n2279);
   U344 : nand3 port map( a => n271, b => n248, c => n268, outb => n270);
   U345 : inv port map( inb => display_out_disp_timer_25_port, outb => n268);
   U346 : aoi12 port map( b => n248, c => display_out_disp_timer_24_port, a => 
                           n272, outb => n269);
   U347 : inv port map( inb => n273, outb => n2280);
   U348 : aoi22 port map( a => n272, b => display_out_disp_timer_24_port, c => 
                           n248, d => n271, outb => n273);
   U349 : inv port map( inb => n274, outb => n272);
   U350 : aoi12 port map( b => n248, c => n275, a => n256, outb => n274);
   U351 : oai22 port map( a => n244, b => n275, c => n276, d => n277, outb => 
                           n2281);
   U352 : aoi12 port map( b => display_out_disp_timer_22_port, c => n248, a => 
                           n278, outb => n276);
   U353 : oai12 port map( b => n279, c => n280, a => n281, outb => n2282);
   U354 : nand3 port map( a => n282, b => n248, c => n280, outb => n281);
   U355 : inv port map( inb => n278, outb => n279);
   U356 : oai12 port map( b => n244, c => n282, a => n265, outb => n278);
   U357 : inv port map( inb => n283, outb => n2283);
   U358 : aoi22 port map( a => n248, b => n282, c => n284, d => 
                           display_out_disp_timer_21_port, outb => n283);
   U359 : oai12 port map( b => n285, c => n244, a => n286, outb => n284);
   U360 : oai12 port map( b => n286, c => n285, a => n287, outb => n2284);
   U361 : nand3 port map( a => n288, b => n248, c => n285, outb => n287);
   U362 : aoi12 port map( b => n248, c => n289, a => n256, outb => n286);
   U363 : inv port map( inb => n290, outb => n2285);
   U364 : aoi22 port map( a => n248, b => n288, c => n291, d => 
                           display_out_disp_timer_19_port, outb => n290);
   U365 : oai12 port map( b => n292, c => n244, a => n293, outb => n291);
   U366 : inv port map( inb => n289, outb => n288);
   U367 : oai12 port map( b => n293, c => n292, a => n294, outb => n2286);
   U368 : nand3 port map( a => n295, b => n248, c => n292, outb => n294);
   U369 : aoi12 port map( b => n248, c => n296, a => n256, outb => n293);
   U370 : oai22 port map( a => n244, b => n296, c => n297, d => n298, outb => 
                           n2287);
   U371 : aoi12 port map( b => display_out_disp_timer_16_port, c => n248, a => 
                           n299, outb => n297);
   U372 : oai12 port map( b => n300, c => n301, a => n302, outb => n2288);
   U373 : nand3 port map( a => n303, b => n248, c => n301, outb => n302);
   U374 : inv port map( inb => n299, outb => n300);
   U375 : oai12 port map( b => n244, c => n303, a => n265, outb => n299);
   U376 : oai12 port map( b => n304, c => n305, a => n306, outb => 
                           load_n_store_n275);
   U377 : aoi22 port map( a => n307, b => n308, c => n309, d => addr_i_0_port, 
                           outb => n306);
   U378 : nor2 port map( a => n310, b => n311, outb => load_n_store_n274);
   U379 : oai12 port map( b => n312, c => n305, a => n313, outb => 
                           load_n_store_n273);
   U380 : aoi22 port map( a => n307, b => n314, c => n309, d => addr_i_4_port, 
                           outb => n313);
   U381 : oai12 port map( b => n315, c => n316, a => n312, outb => n314);
   U382 : inv port map( inb => n317, outb => n316);
   U383 : oai22 port map( a => n318, b => n319, c => n320, d => n321, outb => 
                           load_n_store_n272);
   U384 : inv port map( inb => n320, outb => n318);
   U385 : aoi12 port map( b => n168, c => n322, a => n323, outb => n320);
   U386 : nor3 port map( a => n324, b => n325, c => n326, outb => n323);
   U387 : inv port map( inb => n166, outb => n168);
   U388 : nand2 port map( a => n327, b => n328, outb => load_n_store_n271);
   U389 : oai22 port map( a => n329, b => n310, c => n330, d => n331, outb => 
                           load_n_store_n270);
   U390 : oai22 port map( a => n332, b => n310, c => n333, d => n331, outb => 
                           load_n_store_n269);
   U391 : oai22 port map( a => n334, b => n310, c => n331, d => n335, outb => 
                           load_n_store_n268);
   U392 : inv port map( inb => n336, outb => n335);
   U393 : nand4 port map( a => n337, b => n338, c => top_dv_i, d => n310, outb 
                           => n331);
   U394 : inv port map( inb => n339, outb => n337);
   U395 : inv port map( inb => load_n_store_mem_timer_2_port, outb => n334);
   U396 : nor2 port map( a => n310, b => n340, outb => load_n_store_n267);
   U397 : oai12 port map( b => n341, c => n325, a => n328, outb => n310);
   U398 : aoi12 port map( b => n338, c => n319, a => n342, outb => n341);
   U399 : inv port map( inb => n343, outb => load_n_store_n266);
   U400 : aoi22 port map( a => n344, b => load_n_store_simple_mem_sm_0_port, c 
                           => n345, d => n327, outb => n343);
   U401 : nand4 port map( a => reset_port, b => n346, c => n347, d => n324, 
                           outb => n345);
   U402 : nand3 port map( a => top_dv_i, b => n348, c => n338, outb => n346);
   U403 : inv port map( inb => n327, outb => n344);
   U404 : nand4 port map( a => reset_port, b => n349, c => n350, d => n321, 
                           outb => n327);
   U405 : nand2 port map( a => top_dv_i, b => n351, outb => n349);
   U406 : oai12 port map( b => n325, c => n347, a => n352, outb => 
                           load_n_store_n265);
   U407 : nand2 port map( a => top_ack_port, b => n353, outb => n352);
   U408 : nand4 port map( a => n338, b => n354, c => reset_port, d => n339, 
                           outb => n353);
   U409 : aoi12 port map( b => n355, c => n356, a => n325, outb => 
                           load_n_store_n264);
   U410 : nand3 port map( a => n347, b => n357, c => load_n_store_we_i, outb =>
                           n356);
   U411 : inv port map( inb => n342, outb => n347);
   U412 : nor2 port map( a => n321, b => n354, outb => n342);
   U413 : nand3 port map( a => top_dv_i, b => n358, c => n338, outb => n355);
   U414 : oai12 port map( b => n359, c => n305, a => n360, outb => 
                           load_n_store_n263);
   U415 : aoi22 port map( a => n307, b => n361, c => n309, d => addr_i_1_port, 
                           outb => n360);
   U416 : inv port map( inb => n333, outb => n361);
   U417 : xor2 port map( a => n362, b => n308, outb => n333);
   U418 : inv port map( inb => n330, outb => n308);
   U419 : oai12 port map( b => n363, c => n305, a => n364, outb => 
                           load_n_store_n262);
   U420 : aoi22 port map( a => n336, b => n307, c => n309, d => addr_i_2_port, 
                           outb => n364);
   U421 : xor2 port map( a => n365, b => n366, outb => n336);
   U422 : oai12 port map( b => n315, c => n305, a => n367, outb => 
                           load_n_store_n261);
   U423 : aoi22 port map( a => n368, b => n307, c => n309, d => addr_i_3_port, 
                           outb => n367);
   U424 : nor2 port map( a => n369, b => top_dv_i, outb => n309);
   U425 : nor3 port map( a => n322, b => n369, c => n321, outb => n307);
   U426 : inv port map( inb => n305, outb => n369);
   U427 : nor2 port map( a => n370, b => n371, outb => n322);
   U428 : xor2 port map( a => load_n_store_s_addr_3_port, b => n317, outb => 
                           n368);
   U429 : nor2 port map( a => n365, b => n366, outb => n317);
   U430 : aoi22 port map( a => n372, b => load_n_store_s_addr_2_port, c => 
                           load_n_store_mem_timer_2_port, d => n338, outb => 
                           n366);
   U431 : nand2 port map( a => n362, b => n330, outb => n365);
   U432 : oai22 port map( a => n321, b => n304, c => n329, d => n350, outb => 
                           n330);
   U433 : inv port map( inb => load_n_store_mem_timer_0_port, outb => n329);
   U434 : oai22 port map( a => n321, b => n359, c => n332, d => n350, outb => 
                           n362);
   U435 : inv port map( inb => load_n_store_mem_timer_1_port, outb => n332);
   U436 : inv port map( inb => n372, outb => n321);
   U437 : nand3 port map( a => n166, b => n142, c => n357, outb => n305);
   U438 : nand3 port map( a => n372, b => reset_port, c => n354, outb => n166);
   U439 : nor2 port map( a => n326, b => load_n_store_mem_full, outb => n354);
   U440 : inv port map( inb => top_dv_i, outb => n326);
   U441 : nor2 port map( a => load_n_store_simple_mem_sm_1_port, b => 
                           load_n_store_simple_mem_sm_0_port, outb => n372);
   U442 : nand3 port map( a => n328, b => n142, c => n373, outb => 
                           load_n_store_n260);
   U443 : nand2 port map( a => n374, b => mem_hub_f, outb => n373);
   U444 : nand2 port map( a => n375, b => n351, outb => n142);
   U445 : nand2 port map( a => n338, b => n375, outb => n328);
   U446 : oai22 port map( a => n240, b => n376, c => n374, d => n377, outb => 
                           load_n_store_n259);
   U447 : inv port map( inb => n376, outb => n374);
   U448 : nand3 port map( a => n357, b => n324, c => reset_port, outb => n376);
   U449 : inv port map( inb => n351, outb => n324);
   U450 : nor2 port map( a => n378, b => load_n_store_simple_mem_sm_0_port, 
                           outb => n351);
   U451 : nand2 port map( a => n338, b => n358, outb => n357);
   U452 : oai12 port map( b => n325, c => n348, a => n377, outb => n358);
   U453 : inv port map( inb => n375, outb => n377);
   U454 : nor2 port map( a => n325, b => top_dv_i, outb => n375);
   U455 : nand2 port map( a => n319, b => n339, outb => n348);
   U456 : nand3 port map( a => n340, b => n311, c => n379, outb => n339);
   U457 : nand3 port map( a => load_n_store_mem_timer_1_port, b => 
                           load_n_store_mem_timer_0_port, c => 
                           load_n_store_mem_timer_2_port, outb => n379);
   U458 : inv port map( inb => load_n_store_mem_timer_4_port, outb => n311);
   U459 : inv port map( inb => load_n_store_mem_timer_3_port, outb => n340);
   U460 : inv port map( inb => load_n_store_mem_full, outb => n319);
   U461 : inv port map( inb => reset_port, outb => n325);
   U462 : inv port map( inb => n350, outb => n338);
   U463 : nand2 port map( a => load_n_store_simple_mem_sm_0_port, b => n378, 
                           outb => n350);
   U464 : inv port map( inb => load_n_store_simple_mem_sm_1_port, outb => n378)
                           ;
   U465 : inv port map( inb => mem_reg_f, outb => n240);
   U466 : oai22 port map( a => n177, b => n380, c => n381, d => n382, outb => 
                           n3181);
   U467 : oai22 port map( a => n175, b => n380, c => n381, d => n383, outb => 
                           n3180);
   U468 : oai22 port map( a => n173, b => n380, c => n381, d => n384, outb => 
                           n3179);
   U469 : oai22 port map( a => n171, b => n380, c => n381, d => n385, outb => 
                           n3178);
   U470 : oai22 port map( a => n169, b => n380, c => n381, d => n386, outb => 
                           n3177);
   U471 : oai22 port map( a => n183, b => n387, c => n388, d => n389, outb => 
                           n3176);
   U472 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_10_7_port, 
                           outb => n389);
   U473 : oai22 port map( a => n181, b => n387, c => n388, d => n390, outb => 
                           n3175);
   U474 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_10_6_port, 
                           outb => n390);
   U475 : oai22 port map( a => n179, b => n387, c => n388, d => n391, outb => 
                           n3174);
   U476 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_10_5_port, 
                           outb => n391);
   U477 : oai22 port map( a => n177, b => n387, c => n388, d => n392, outb => 
                           n3173);
   U478 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_10_4_port, 
                           outb => n392);
   U479 : oai22 port map( a => n175, b => n387, c => n388, d => n393, outb => 
                           n3172);
   U480 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_10_3_port, 
                           outb => n393);
   U481 : oai22 port map( a => n173, b => n387, c => n388, d => n394, outb => 
                           n3171);
   U482 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_10_2_port, 
                           outb => n394);
   U483 : oai22 port map( a => n171, b => n387, c => n388, d => n395, outb => 
                           n3170);
   U484 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_10_1_port, 
                           outb => n395);
   U485 : oai22 port map( a => n169, b => n387, c => n388, d => n396, outb => 
                           n3169);
   U486 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_10_0_port, 
                           outb => n396);
   U487 : oai22 port map( a => n183, b => n397, c => n398, d => n399, outb => 
                           n3168);
   U488 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_9_7_port, 
                           outb => n399);
   U489 : oai22 port map( a => n181, b => n397, c => n398, d => n400, outb => 
                           n3167);
   U490 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_9_6_port, 
                           outb => n400);
   U491 : oai22 port map( a => n179, b => n397, c => n398, d => n401, outb => 
                           n3166);
   U492 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_9_5_port, 
                           outb => n401);
   U493 : oai22 port map( a => n177, b => n397, c => n398, d => n402, outb => 
                           n3165);
   U494 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_9_4_port, 
                           outb => n402);
   U495 : oai22 port map( a => n175, b => n397, c => n398, d => n403, outb => 
                           n3164);
   U496 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_9_3_port, 
                           outb => n403);
   U497 : oai22 port map( a => n173, b => n397, c => n398, d => n404, outb => 
                           n3163);
   U498 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_9_2_port, 
                           outb => n404);
   U499 : oai22 port map( a => n171, b => n397, c => n398, d => n405, outb => 
                           n3162);
   U500 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_9_1_port, 
                           outb => n405);
   U501 : oai22 port map( a => n169, b => n397, c => n398, d => n406, outb => 
                           n3161);
   U502 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_9_0_port, 
                           outb => n406);
   U503 : oai22 port map( a => n183, b => n407, c => n408, d => n409, outb => 
                           n3160);
   U504 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_8_7_port, 
                           outb => n409);
   U505 : oai22 port map( a => n181, b => n407, c => n408, d => n410, outb => 
                           n3159);
   U506 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_8_6_port, 
                           outb => n410);
   U507 : oai22 port map( a => n179, b => n407, c => n408, d => n411, outb => 
                           n3158);
   U508 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_8_5_port, 
                           outb => n411);
   U509 : oai22 port map( a => n177, b => n407, c => n408, d => n412, outb => 
                           n3157);
   U510 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_8_4_port, 
                           outb => n412);
   U511 : oai22 port map( a => n175, b => n407, c => n408, d => n413, outb => 
                           n3156);
   U512 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_8_3_port, 
                           outb => n413);
   U513 : oai22 port map( a => n173, b => n407, c => n408, d => n414, outb => 
                           n3155);
   U514 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_8_2_port, 
                           outb => n414);
   U515 : oai22 port map( a => n171, b => n407, c => n408, d => n415, outb => 
                           n3154);
   U516 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_8_1_port, 
                           outb => n415);
   U517 : oai22 port map( a => n169, b => n407, c => n408, d => n416, outb => 
                           n3153);
   U518 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_8_0_port, 
                           outb => n416);
   U519 : oai22 port map( a => n183, b => n417, c => n418, d => n419, outb => 
                           n3152);
   U520 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_7_7_port, 
                           outb => n419);
   U521 : oai22 port map( a => n181, b => n417, c => n418, d => n420, outb => 
                           n3151);
   U522 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_7_6_port, 
                           outb => n420);
   U523 : oai22 port map( a => n179, b => n417, c => n418, d => n421, outb => 
                           n3150);
   U524 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_7_5_port, 
                           outb => n421);
   U525 : oai22 port map( a => n177, b => n417, c => n418, d => n422, outb => 
                           n3149);
   U526 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_7_4_port, 
                           outb => n422);
   U527 : oai22 port map( a => n175, b => n417, c => n418, d => n423, outb => 
                           n3148);
   U528 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_7_3_port, 
                           outb => n423);
   U529 : oai22 port map( a => n173, b => n417, c => n418, d => n424, outb => 
                           n3147);
   U530 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_7_2_port, 
                           outb => n424);
   U531 : oai22 port map( a => n171, b => n417, c => n418, d => n425, outb => 
                           n3146);
   U532 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_7_1_port, 
                           outb => n425);
   U533 : oai22 port map( a => n169, b => n417, c => n418, d => n426, outb => 
                           n3145);
   U534 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_7_0_port, 
                           outb => n426);
   U535 : oai22 port map( a => n183, b => n427, c => n428, d => n429, outb => 
                           n3144);
   U536 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_6_7_port, 
                           outb => n429);
   U537 : oai22 port map( a => n181, b => n427, c => n428, d => n430, outb => 
                           n3143);
   U538 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_6_6_port, 
                           outb => n430);
   U539 : oai22 port map( a => n179, b => n427, c => n428, d => n431, outb => 
                           n3142);
   U540 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_6_5_port, 
                           outb => n431);
   U541 : oai22 port map( a => n177, b => n427, c => n428, d => n432, outb => 
                           n3141);
   U542 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_6_4_port, 
                           outb => n432);
   U543 : oai22 port map( a => n175, b => n427, c => n428, d => n433, outb => 
                           n3140);
   U544 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_6_3_port, 
                           outb => n433);
   U545 : oai22 port map( a => n173, b => n427, c => n428, d => n434, outb => 
                           n3139);
   U546 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_6_2_port, 
                           outb => n434);
   U547 : oai22 port map( a => n171, b => n427, c => n428, d => n435, outb => 
                           n3138);
   U548 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_6_1_port, 
                           outb => n435);
   U549 : oai22 port map( a => n169, b => n427, c => n428, d => n436, outb => 
                           n3137);
   U550 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_6_0_port, 
                           outb => n436);
   U551 : oai22 port map( a => n183, b => n437, c => n438, d => n439, outb => 
                           n3136);
   U552 : oai22 port map( a => n181, b => n437, c => n438, d => n440, outb => 
                           n3135);
   U553 : oai22 port map( a => n179, b => n437, c => n438, d => n441, outb => 
                           n3134);
   U554 : oai22 port map( a => n177, b => n437, c => n438, d => n442, outb => 
                           n3133);
   U555 : oai22 port map( a => n175, b => n437, c => n438, d => n443, outb => 
                           n3132);
   U556 : oai22 port map( a => n173, b => n437, c => n438, d => n444, outb => 
                           n3131);
   U557 : oai22 port map( a => n171, b => n437, c => n438, d => n445, outb => 
                           n3130);
   U558 : oai22 port map( a => n169, b => n437, c => n438, d => n446, outb => 
                           n3129);
   U559 : oai22 port map( a => n183, b => n447, c => n448, d => n449, outb => 
                           n3128);
   U560 : oai22 port map( a => n181, b => n447, c => n448, d => n450, outb => 
                           n3127);
   U561 : oai22 port map( a => n179, b => n447, c => n448, d => n451, outb => 
                           n3126);
   U562 : oai22 port map( a => n177, b => n447, c => n448, d => n452, outb => 
                           n3125);
   U563 : oai22 port map( a => n175, b => n447, c => n448, d => n453, outb => 
                           n3124);
   U564 : oai22 port map( a => n173, b => n447, c => n448, d => n454, outb => 
                           n3123);
   U565 : oai22 port map( a => n171, b => n447, c => n448, d => n455, outb => 
                           n3122);
   U566 : oai22 port map( a => n169, b => n447, c => n448, d => n456, outb => 
                           n3121);
   U567 : oai22 port map( a => n183, b => n457, c => n458, d => n459, outb => 
                           n3120);
   U568 : oai22 port map( a => n181, b => n457, c => n458, d => n460, outb => 
                           n3119);
   U569 : oai22 port map( a => n179, b => n457, c => n458, d => n461, outb => 
                           n3118);
   U570 : oai22 port map( a => n177, b => n457, c => n458, d => n462, outb => 
                           n3117);
   U571 : oai22 port map( a => n175, b => n457, c => n458, d => n463, outb => 
                           n3116);
   U572 : oai22 port map( a => n173, b => n457, c => n458, d => n464, outb => 
                           n3115);
   U573 : oai22 port map( a => n171, b => n457, c => n458, d => n465, outb => 
                           n3114);
   U574 : oai22 port map( a => n169, b => n457, c => n458, d => n466, outb => 
                           n3113);
   U575 : oai22 port map( a => n183, b => n467, c => n468, d => n469, outb => 
                           n3112);
   U576 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_2_7_port, 
                           outb => n469);
   U577 : oai22 port map( a => n181, b => n467, c => n468, d => n470, outb => 
                           n3111);
   U578 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_2_6_port, 
                           outb => n470);
   U579 : oai22 port map( a => n179, b => n467, c => n468, d => n471, outb => 
                           n3110);
   U580 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_2_5_port, 
                           outb => n471);
   U581 : oai22 port map( a => n177, b => n467, c => n468, d => n472, outb => 
                           n3109);
   U582 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_2_4_port, 
                           outb => n472);
   U583 : oai22 port map( a => n175, b => n467, c => n468, d => n473, outb => 
                           n3108);
   U584 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_2_3_port, 
                           outb => n473);
   U585 : oai22 port map( a => n173, b => n467, c => n468, d => n474, outb => 
                           n3107);
   U586 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_2_2_port, 
                           outb => n474);
   U587 : oai22 port map( a => n171, b => n467, c => n468, d => n475, outb => 
                           n3106);
   U588 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_2_1_port, 
                           outb => n475);
   U589 : oai22 port map( a => n169, b => n467, c => n468, d => n476, outb => 
                           n3105);
   U590 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_2_0_port, 
                           outb => n476);
   U591 : oai22 port map( a => n183, b => n477, c => n478, d => n479, outb => 
                           n3104);
   U592 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_1_7_port, 
                           outb => n479);
   U593 : oai22 port map( a => n181, b => n477, c => n478, d => n480, outb => 
                           n3103);
   U594 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_1_6_port, 
                           outb => n480);
   U595 : oai22 port map( a => n179, b => n477, c => n478, d => n481, outb => 
                           n3102);
   U596 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_1_5_port, 
                           outb => n481);
   U597 : oai22 port map( a => n177, b => n477, c => n478, d => n482, outb => 
                           n3101);
   U598 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_1_4_port, 
                           outb => n482);
   U599 : oai22 port map( a => n175, b => n477, c => n478, d => n483, outb => 
                           n3100);
   U600 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_1_3_port, 
                           outb => n483);
   U601 : oai22 port map( a => n173, b => n477, c => n478, d => n484, outb => 
                           n3099);
   U602 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_1_2_port, 
                           outb => n484);
   U603 : oai22 port map( a => n171, b => n477, c => n478, d => n485, outb => 
                           n3098);
   U604 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_1_1_port, 
                           outb => n485);
   U605 : oai22 port map( a => n169, b => n477, c => n478, d => n486, outb => 
                           n3097);
   U606 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_1_0_port, 
                           outb => n486);
   U607 : oai22 port map( a => n183, b => n487, c => n488, d => n489, outb => 
                           n3096);
   U608 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_0_7_port, 
                           outb => n489);
   U609 : oai22 port map( a => n181, b => n487, c => n488, d => n490, outb => 
                           n3095);
   U610 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_0_6_port, 
                           outb => n490);
   U611 : oai22 port map( a => n179, b => n487, c => n488, d => n491, outb => 
                           n3094);
   U612 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_0_5_port, 
                           outb => n491);
   U613 : oai22 port map( a => n177, b => n487, c => n488, d => n492, outb => 
                           n3093);
   U614 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_0_4_port, 
                           outb => n492);
   U615 : oai22 port map( a => n175, b => n487, c => n488, d => n493, outb => 
                           n3092);
   U616 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_0_3_port, 
                           outb => n493);
   U617 : oai22 port map( a => n173, b => n487, c => n488, d => n494, outb => 
                           n3091);
   U618 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_0_2_port, 
                           outb => n494);
   U619 : oai22 port map( a => n171, b => n487, c => n488, d => n495, outb => 
                           n3090);
   U620 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_0_1_port, 
                           outb => n495);
   U621 : oai22 port map( a => n169, b => n487, c => n488, d => n496, outb => 
                           n3089);
   U622 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_0_0_port, 
                           outb => n496);
   U623 : nand4 port map( a => n497, b => n498, c => n499, d => n500, outb => 
                           n2839);
   U624 : aoi22 port map( a => n501, b => n502, c => load_n_store_we_i, d => 
                           load_n_store_lazy_in_2_7_port, outb => n500);
   U625 : nor3 port map( a => n503, b => n504, c => n505, outb => n502);
   U626 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_26_7_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_31_7_port, d =>
                           n370, outb => n505);
   U627 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_25_7_port, b
                           => n507, outb => n504);
   U628 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_30_7_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_24_7_port, d =>
                           n509, outb => n503);
   U629 : nor3 port map( a => n510, b => n511, c => n512, outb => n501);
   U630 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_27_7_port, b
                           => n513, outb => n511);
   U631 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_28_7_port, 
                           b => n514, c => 
                           load_n_store_RGB_Array_2_block_ram_r_29_7_port, d =>
                           n515, outb => n510);
   U632 : nand4 port map( a => n516, b => n517, c => n518, d => n519, outb => 
                           n499);
   U633 : nor3 port map( a => n520, b => n521, c => n522, outb => n519);
   U634 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_18_7_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_23_7_port, d =>
                           n370, outb => n522);
   U635 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_17_7_port, b
                           => n507, outb => n521);
   U636 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_22_7_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_16_7_port, d =>
                           n509, outb => n520);
   U637 : aoi22 port map( a => n523, b => n524, c => n525, d => n526, outb => 
                           n518);
   U638 : nand2 port map( a => n527, b => n528, outb => n517);
   U639 : nand4 port map( a => n529, b => n530, c => n531, d => n532, outb => 
                           n498);
   U640 : nor3 port map( a => n533, b => n534, c => n535, outb => n532);
   U641 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_10_7_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_15_7_port, d =>
                           n370, outb => n535);
   U642 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_9_7_port, b 
                           => n507, outb => n534);
   U643 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_14_7_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_8_7_port, d => 
                           n509, outb => n533);
   U644 : aoi22 port map( a => n523, b => n536, c => n525, d => n537, outb => 
                           n531);
   U645 : nand2 port map( a => n527, b => n538, outb => n530);
   U646 : nand4 port map( a => n539, b => n540, c => n541, d => n542, outb => 
                           n497);
   U647 : nor3 port map( a => n543, b => n544, c => n545, outb => n542);
   U648 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_2_7_port, b
                           => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_7_7_port, d => 
                           n370, outb => n545);
   U649 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_1_7_port, b 
                           => n507, outb => n544);
   U650 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_6_7_port, b
                           => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_0_7_port, d => 
                           n509, outb => n543);
   U651 : aoi22 port map( a => n523, b => n439, c => n525, d => n449, outb => 
                           n541);
   U652 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_4_7_port, 
                           outb => n449);
   U653 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_5_7_port, 
                           outb => n439);
   U654 : nand2 port map( a => n527, b => n459, outb => n540);
   U655 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_3_7_port, 
                           outb => n459);
   U656 : nand4 port map( a => n546, b => n547, c => n548, d => n549, outb => 
                           n2836);
   U657 : aoi22 port map( a => n550, b => n551, c => load_n_store_we_i, d => 
                           load_n_store_lazy_in_2_6_port, outb => n549);
   U658 : nor3 port map( a => n552, b => n553, c => n554, outb => n551);
   U659 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_26_6_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_31_6_port, d =>
                           n370, outb => n554);
   U660 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_25_6_port, b
                           => n507, outb => n553);
   U661 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_30_6_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_24_6_port, d =>
                           n509, outb => n552);
   U662 : nor3 port map( a => n555, b => n556, c => n512, outb => n550);
   U663 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_27_6_port, b
                           => n513, outb => n556);
   U664 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_28_6_port, 
                           b => n514, c => 
                           load_n_store_RGB_Array_2_block_ram_r_29_6_port, d =>
                           n515, outb => n555);
   U665 : nand4 port map( a => n516, b => n557, c => n558, d => n559, outb => 
                           n548);
   U666 : nor3 port map( a => n560, b => n561, c => n562, outb => n559);
   U667 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_18_6_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_23_6_port, d =>
                           n370, outb => n562);
   U668 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_17_6_port, b
                           => n507, outb => n561);
   U669 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_22_6_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_16_6_port, d =>
                           n509, outb => n560);
   U670 : aoi22 port map( a => n523, b => n563, c => n525, d => n564, outb => 
                           n558);
   U671 : nand2 port map( a => n527, b => n565, outb => n557);
   U672 : nand4 port map( a => n529, b => n566, c => n567, d => n568, outb => 
                           n547);
   U673 : nor3 port map( a => n569, b => n570, c => n571, outb => n568);
   U674 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_10_6_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_15_6_port, d =>
                           n370, outb => n571);
   U675 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_9_6_port, b 
                           => n507, outb => n570);
   U676 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_14_6_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_8_6_port, d => 
                           n509, outb => n569);
   U677 : aoi22 port map( a => n523, b => n572, c => n525, d => n573, outb => 
                           n567);
   U678 : nand2 port map( a => n527, b => n574, outb => n566);
   U679 : nand4 port map( a => n539, b => n575, c => n576, d => n577, outb => 
                           n546);
   U680 : nor3 port map( a => n578, b => n579, c => n580, outb => n577);
   U681 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_2_6_port, b
                           => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_7_6_port, d => 
                           n370, outb => n580);
   U682 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_1_6_port, b 
                           => n507, outb => n579);
   U683 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_6_6_port, b
                           => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_0_6_port, d => 
                           n509, outb => n578);
   U684 : aoi22 port map( a => n523, b => n440, c => n525, d => n450, outb => 
                           n576);
   U685 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_4_6_port, 
                           outb => n450);
   U686 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_5_6_port, 
                           outb => n440);
   U687 : nand2 port map( a => n527, b => n460, outb => n575);
   U688 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_3_6_port, 
                           outb => n460);
   U689 : nand4 port map( a => n581, b => n582, c => n583, d => n584, outb => 
                           n2833);
   U690 : aoi22 port map( a => n585, b => n586, c => load_n_store_we_i, d => 
                           load_n_store_lazy_in_2_5_port, outb => n584);
   U691 : nor3 port map( a => n587, b => n588, c => n589, outb => n586);
   U692 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_26_5_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_31_5_port, d =>
                           n370, outb => n589);
   U693 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_25_5_port, b
                           => n507, outb => n588);
   U694 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_30_5_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_24_5_port, d =>
                           n509, outb => n587);
   U695 : nor3 port map( a => n590, b => n591, c => n512, outb => n585);
   U696 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_27_5_port, b
                           => n513, outb => n591);
   U697 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_28_5_port, 
                           b => n514, c => 
                           load_n_store_RGB_Array_2_block_ram_r_29_5_port, d =>
                           n515, outb => n590);
   U698 : nand4 port map( a => n516, b => n592, c => n593, d => n594, outb => 
                           n583);
   U699 : nor3 port map( a => n595, b => n596, c => n597, outb => n594);
   U700 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_18_5_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_23_5_port, d =>
                           n370, outb => n597);
   U701 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_17_5_port, b
                           => n507, outb => n596);
   U702 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_22_5_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_16_5_port, d =>
                           n509, outb => n595);
   U703 : aoi22 port map( a => n523, b => n598, c => n525, d => n599, outb => 
                           n593);
   U704 : nand2 port map( a => n527, b => n600, outb => n592);
   U705 : nand4 port map( a => n529, b => n601, c => n602, d => n603, outb => 
                           n582);
   U706 : nor3 port map( a => n604, b => n605, c => n606, outb => n603);
   U707 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_10_5_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_15_5_port, d =>
                           n370, outb => n606);
   U708 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_9_5_port, b 
                           => n507, outb => n605);
   U709 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_14_5_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_8_5_port, d => 
                           n509, outb => n604);
   U710 : aoi22 port map( a => n523, b => n607, c => n525, d => n608, outb => 
                           n602);
   U711 : nand2 port map( a => n527, b => n609, outb => n601);
   U712 : nand4 port map( a => n539, b => n610, c => n611, d => n612, outb => 
                           n581);
   U713 : nor3 port map( a => n613, b => n614, c => n615, outb => n612);
   U714 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_2_5_port, b
                           => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_7_5_port, d => 
                           n370, outb => n615);
   U715 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_1_5_port, b 
                           => n507, outb => n614);
   U716 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_6_5_port, b
                           => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_0_5_port, d => 
                           n509, outb => n613);
   U717 : aoi22 port map( a => n523, b => n441, c => n525, d => n451, outb => 
                           n611);
   U718 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_4_5_port, 
                           outb => n451);
   U719 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_5_5_port, 
                           outb => n441);
   U720 : nand2 port map( a => n527, b => n461, outb => n610);
   U721 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_3_5_port, 
                           outb => n461);
   U722 : nand4 port map( a => n616, b => n617, c => n618, d => n619, outb => 
                           n2830);
   U723 : aoi22 port map( a => n620, b => n621, c => load_n_store_we_i, d => 
                           load_n_store_lazy_in_2_4_port, outb => n619);
   U724 : nor3 port map( a => n622, b => n623, c => n624, outb => n621);
   U725 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_26_4_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_31_4_port, d =>
                           n370, outb => n624);
   U726 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_25_4_port, b
                           => n507, outb => n623);
   U727 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_30_4_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_24_4_port, d =>
                           n509, outb => n622);
   U728 : nor3 port map( a => n625, b => n626, c => n512, outb => n620);
   U729 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_27_4_port, b
                           => n513, outb => n626);
   U730 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_28_4_port, 
                           b => n514, c => 
                           load_n_store_RGB_Array_2_block_ram_r_29_4_port, d =>
                           n515, outb => n625);
   U731 : nand4 port map( a => n516, b => n627, c => n628, d => n629, outb => 
                           n618);
   U732 : nor3 port map( a => n630, b => n631, c => n632, outb => n629);
   U733 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_18_4_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_23_4_port, d =>
                           n370, outb => n632);
   U734 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_17_4_port, b
                           => n507, outb => n631);
   U735 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_22_4_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_16_4_port, d =>
                           n509, outb => n630);
   U736 : aoi22 port map( a => n523, b => n633, c => n525, d => n634, outb => 
                           n628);
   U737 : nand2 port map( a => n527, b => n635, outb => n627);
   U738 : nand4 port map( a => n529, b => n636, c => n637, d => n638, outb => 
                           n617);
   U739 : nor3 port map( a => n639, b => n640, c => n641, outb => n638);
   U740 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_10_4_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_15_4_port, d =>
                           n370, outb => n641);
   U741 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_9_4_port, b 
                           => n507, outb => n640);
   U742 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_14_4_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_8_4_port, d => 
                           n509, outb => n639);
   U743 : aoi22 port map( a => n523, b => n642, c => n525, d => n643, outb => 
                           n637);
   U744 : nand2 port map( a => n527, b => n382, outb => n636);
   U745 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_11_4_port, 
                           outb => n382);
   U746 : nand4 port map( a => n539, b => n644, c => n645, d => n646, outb => 
                           n616);
   U747 : nor3 port map( a => n647, b => n648, c => n649, outb => n646);
   U748 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_2_4_port, b
                           => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_7_4_port, d => 
                           n370, outb => n649);
   U749 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_1_4_port, b 
                           => n507, outb => n648);
   U750 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_6_4_port, b
                           => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_0_4_port, d => 
                           n509, outb => n647);
   U751 : aoi22 port map( a => n523, b => n442, c => n525, d => n452, outb => 
                           n645);
   U752 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_4_4_port, 
                           outb => n452);
   U753 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_5_4_port, 
                           outb => n442);
   U754 : nand2 port map( a => n527, b => n462, outb => n644);
   U755 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_3_4_port, 
                           outb => n462);
   U756 : nand4 port map( a => n650, b => n651, c => n652, d => n653, outb => 
                           n2827);
   U757 : aoi22 port map( a => n654, b => n655, c => load_n_store_we_i, d => 
                           load_n_store_lazy_in_2_3_port, outb => n653);
   U758 : nor3 port map( a => n656, b => n657, c => n658, outb => n655);
   U759 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_26_3_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_31_3_port, d =>
                           n370, outb => n658);
   U760 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_25_3_port, b
                           => n507, outb => n657);
   U761 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_30_3_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_24_3_port, d =>
                           n509, outb => n656);
   U762 : nor3 port map( a => n659, b => n660, c => n512, outb => n654);
   U763 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_27_3_port, b
                           => n513, outb => n660);
   U764 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_28_3_port, 
                           b => n514, c => 
                           load_n_store_RGB_Array_2_block_ram_r_29_3_port, d =>
                           n515, outb => n659);
   U765 : nand4 port map( a => n516, b => n661, c => n662, d => n663, outb => 
                           n652);
   U766 : nor3 port map( a => n664, b => n665, c => n666, outb => n663);
   U767 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_18_3_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_23_3_port, d =>
                           n370, outb => n666);
   U768 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_17_3_port, b
                           => n507, outb => n665);
   U769 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_22_3_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_16_3_port, d =>
                           n509, outb => n664);
   U770 : aoi22 port map( a => n523, b => n667, c => n525, d => n668, outb => 
                           n662);
   U771 : nand2 port map( a => n527, b => n669, outb => n661);
   U772 : nand4 port map( a => n529, b => n670, c => n671, d => n672, outb => 
                           n651);
   U773 : nor3 port map( a => n673, b => n674, c => n675, outb => n672);
   U774 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_10_3_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_15_3_port, d =>
                           n370, outb => n675);
   U775 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_9_3_port, b 
                           => n507, outb => n674);
   U776 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_14_3_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_8_3_port, d => 
                           n509, outb => n673);
   U777 : aoi22 port map( a => n523, b => n676, c => n525, d => n677, outb => 
                           n671);
   U778 : nand2 port map( a => n527, b => n383, outb => n670);
   U779 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_11_3_port, 
                           outb => n383);
   U780 : nand4 port map( a => n539, b => n678, c => n679, d => n680, outb => 
                           n650);
   U781 : nor3 port map( a => n681, b => n682, c => n683, outb => n680);
   U782 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_2_3_port, b
                           => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_7_3_port, d => 
                           n370, outb => n683);
   U783 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_1_3_port, b 
                           => n507, outb => n682);
   U784 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_6_3_port, b
                           => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_0_3_port, d => 
                           n509, outb => n681);
   U785 : aoi22 port map( a => n523, b => n443, c => n525, d => n453, outb => 
                           n679);
   U786 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_4_3_port, 
                           outb => n453);
   U787 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_5_3_port, 
                           outb => n443);
   U788 : nand2 port map( a => n527, b => n463, outb => n678);
   U789 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_3_3_port, 
                           outb => n463);
   U790 : nand4 port map( a => n684, b => n685, c => n686, d => n687, outb => 
                           n2824);
   U791 : aoi22 port map( a => n688, b => n689, c => load_n_store_we_i, d => 
                           load_n_store_lazy_in_2_2_port, outb => n687);
   U792 : nor3 port map( a => n690, b => n691, c => n692, outb => n689);
   U793 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_26_2_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_31_2_port, d =>
                           n370, outb => n692);
   U794 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_25_2_port, b
                           => n507, outb => n691);
   U795 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_30_2_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_24_2_port, d =>
                           n509, outb => n690);
   U796 : nor3 port map( a => n693, b => n694, c => n512, outb => n688);
   U797 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_27_2_port, b
                           => n513, outb => n694);
   U798 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_28_2_port, 
                           b => n514, c => 
                           load_n_store_RGB_Array_2_block_ram_r_29_2_port, d =>
                           n515, outb => n693);
   U799 : nand4 port map( a => n516, b => n695, c => n696, d => n697, outb => 
                           n686);
   U800 : nor3 port map( a => n698, b => n699, c => n700, outb => n697);
   U801 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_18_2_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_23_2_port, d =>
                           n370, outb => n700);
   U802 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_17_2_port, b
                           => n507, outb => n699);
   U803 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_22_2_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_16_2_port, d =>
                           n509, outb => n698);
   U804 : aoi22 port map( a => n523, b => n701, c => n525, d => n702, outb => 
                           n696);
   U805 : nand2 port map( a => n527, b => n703, outb => n695);
   U806 : nand4 port map( a => n529, b => n704, c => n705, d => n706, outb => 
                           n685);
   U807 : nor3 port map( a => n707, b => n708, c => n709, outb => n706);
   U808 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_10_2_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_15_2_port, d =>
                           n370, outb => n709);
   U809 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_9_2_port, b 
                           => n507, outb => n708);
   U810 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_14_2_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_8_2_port, d => 
                           n509, outb => n707);
   U811 : aoi22 port map( a => n523, b => n710, c => n525, d => n711, outb => 
                           n705);
   U812 : nand2 port map( a => n527, b => n384, outb => n704);
   U813 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_11_2_port, 
                           outb => n384);
   U814 : nand4 port map( a => n539, b => n712, c => n713, d => n714, outb => 
                           n684);
   U815 : nor3 port map( a => n715, b => n716, c => n717, outb => n714);
   U816 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_2_2_port, b
                           => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_7_2_port, d => 
                           n370, outb => n717);
   U817 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_1_2_port, b 
                           => n507, outb => n716);
   U818 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_6_2_port, b
                           => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_0_2_port, d => 
                           n509, outb => n715);
   U819 : aoi22 port map( a => n523, b => n444, c => n525, d => n454, outb => 
                           n713);
   U820 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_4_2_port, 
                           outb => n454);
   U821 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_5_2_port, 
                           outb => n444);
   U822 : nand2 port map( a => n527, b => n464, outb => n712);
   U823 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_3_2_port, 
                           outb => n464);
   U824 : nand4 port map( a => n718, b => n719, c => n720, d => n721, outb => 
                           n2821);
   U825 : aoi22 port map( a => n722, b => n723, c => load_n_store_we_i, d => 
                           load_n_store_lazy_in_2_1_port, outb => n721);
   U826 : nor3 port map( a => n724, b => n725, c => n726, outb => n723);
   U827 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_26_1_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_31_1_port, d =>
                           n370, outb => n726);
   U828 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_25_1_port, b
                           => n507, outb => n725);
   U829 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_30_1_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_24_1_port, d =>
                           n509, outb => n724);
   U830 : nor3 port map( a => n727, b => n728, c => n512, outb => n722);
   U831 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_27_1_port, b
                           => n513, outb => n728);
   U832 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_28_1_port, 
                           b => n514, c => 
                           load_n_store_RGB_Array_2_block_ram_r_29_1_port, d =>
                           n515, outb => n727);
   U833 : nand4 port map( a => n516, b => n729, c => n730, d => n731, outb => 
                           n720);
   U834 : nor3 port map( a => n732, b => n733, c => n734, outb => n731);
   U835 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_18_1_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_23_1_port, d =>
                           n370, outb => n734);
   U836 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_17_1_port, b
                           => n507, outb => n733);
   U837 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_22_1_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_16_1_port, d =>
                           n509, outb => n732);
   U838 : aoi22 port map( a => n523, b => n735, c => n525, d => n736, outb => 
                           n730);
   U839 : nand2 port map( a => n527, b => n737, outb => n729);
   U840 : nand4 port map( a => n529, b => n738, c => n739, d => n740, outb => 
                           n719);
   U841 : nor3 port map( a => n741, b => n742, c => n743, outb => n740);
   U842 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_10_1_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_15_1_port, d =>
                           n370, outb => n743);
   U843 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_9_1_port, b 
                           => n507, outb => n742);
   U844 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_14_1_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_8_1_port, d => 
                           n509, outb => n741);
   U845 : aoi22 port map( a => n523, b => n744, c => n525, d => n745, outb => 
                           n739);
   U846 : nand2 port map( a => n527, b => n385, outb => n738);
   U847 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_11_1_port, 
                           outb => n385);
   U848 : nand4 port map( a => n539, b => n746, c => n747, d => n748, outb => 
                           n718);
   U849 : nor3 port map( a => n749, b => n750, c => n751, outb => n748);
   U850 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_2_1_port, b
                           => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_7_1_port, d => 
                           n370, outb => n751);
   U851 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_1_1_port, b 
                           => n507, outb => n750);
   U852 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_6_1_port, b
                           => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_0_1_port, d => 
                           n509, outb => n749);
   U853 : aoi22 port map( a => n523, b => n445, c => n525, d => n455, outb => 
                           n747);
   U854 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_4_1_port, 
                           outb => n455);
   U855 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_5_1_port, 
                           outb => n445);
   U856 : nand2 port map( a => n527, b => n465, outb => n746);
   U857 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_3_1_port, 
                           outb => n465);
   U858 : nand4 port map( a => n752, b => n753, c => n754, d => n755, outb => 
                           n2818);
   U859 : aoi22 port map( a => n756, b => n757, c => load_n_store_we_i, d => 
                           load_n_store_lazy_in_2_0_port, outb => n755);
   U860 : nor3 port map( a => n758, b => n759, c => n760, outb => n757);
   U861 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_26_0_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_31_0_port, d =>
                           n370, outb => n760);
   U862 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_25_0_port, b
                           => n507, outb => n759);
   U863 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_30_0_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_24_0_port, d =>
                           n509, outb => n758);
   U864 : nor3 port map( a => n761, b => n762, c => n512, outb => n756);
   U865 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_27_0_port, b
                           => n513, outb => n762);
   U866 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_28_0_port, 
                           b => n514, c => 
                           load_n_store_RGB_Array_2_block_ram_r_29_0_port, d =>
                           n515, outb => n761);
   U867 : nand4 port map( a => n516, b => n763, c => n764, d => n765, outb => 
                           n754);
   U868 : nor3 port map( a => n766, b => n767, c => n768, outb => n765);
   U869 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_18_0_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_23_0_port, d =>
                           n370, outb => n768);
   U870 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_17_0_port, b
                           => n507, outb => n767);
   U871 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_22_0_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_16_0_port, d =>
                           n509, outb => n766);
   U872 : aoi22 port map( a => n523, b => n769, c => n525, d => n770, outb => 
                           n764);
   U873 : nand2 port map( a => n527, b => n771, outb => n763);
   U874 : nand4 port map( a => n529, b => n772, c => n773, d => n774, outb => 
                           n753);
   U875 : nor3 port map( a => n775, b => n776, c => n777, outb => n774);
   U876 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_10_0_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_15_0_port, d =>
                           n370, outb => n777);
   U877 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_9_0_port, b 
                           => n507, outb => n776);
   U878 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_14_0_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_8_0_port, d => 
                           n509, outb => n775);
   U879 : aoi22 port map( a => n523, b => n778, c => n525, d => n779, outb => 
                           n773);
   U880 : nand2 port map( a => n527, b => n386, outb => n772);
   U881 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_11_0_port, 
                           outb => n386);
   U882 : nand4 port map( a => n539, b => n780, c => n781, d => n782, outb => 
                           n752);
   U883 : nor3 port map( a => n783, b => n784, c => n785, outb => n782);
   U884 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_2_0_port, b
                           => n506, c => 
                           load_n_store_RGB_Array_2_block_ram_r_7_0_port, d => 
                           n370, outb => n785);
   U885 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_1_0_port, b 
                           => n507, outb => n784);
   U886 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_6_0_port, b
                           => n508, c => 
                           load_n_store_RGB_Array_2_block_ram_r_0_0_port, d => 
                           n509, outb => n783);
   U887 : aoi22 port map( a => n523, b => n446, c => n525, d => n456, outb => 
                           n781);
   U888 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_4_0_port, 
                           outb => n456);
   U889 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_5_0_port, 
                           outb => n446);
   U890 : nand2 port map( a => n527, b => n466, outb => n780);
   U891 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_3_0_port, 
                           outb => n466);
   U892 : oai22 port map( a => n183, b => n786, c => n787, d => n788, outb => 
                           n3344);
   U893 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_31_7_port, 
                           outb => n788);
   U894 : oai22 port map( a => n181, b => n786, c => n787, d => n789, outb => 
                           n3343);
   U895 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_31_6_port, 
                           outb => n789);
   U896 : oai22 port map( a => n179, b => n786, c => n787, d => n790, outb => 
                           n3342);
   U897 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_31_5_port, 
                           outb => n790);
   U898 : oai22 port map( a => n177, b => n786, c => n787, d => n791, outb => 
                           n3341);
   U899 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_31_4_port, 
                           outb => n791);
   U900 : oai22 port map( a => n175, b => n786, c => n787, d => n792, outb => 
                           n3340);
   U901 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_31_3_port, 
                           outb => n792);
   U902 : oai22 port map( a => n173, b => n786, c => n787, d => n793, outb => 
                           n3339);
   U903 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_31_2_port, 
                           outb => n793);
   U904 : oai22 port map( a => n171, b => n786, c => n787, d => n794, outb => 
                           n3338);
   U905 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_31_1_port, 
                           outb => n794);
   U906 : oai22 port map( a => n169, b => n786, c => n787, d => n795, outb => 
                           n3337);
   U907 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_31_0_port, 
                           outb => n795);
   U908 : oai22 port map( a => n183, b => n796, c => n797, d => n798, outb => 
                           n3336);
   U909 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_30_7_port, 
                           outb => n798);
   U910 : oai22 port map( a => n181, b => n796, c => n797, d => n799, outb => 
                           n3335);
   U911 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_30_6_port, 
                           outb => n799);
   U912 : oai22 port map( a => n179, b => n796, c => n797, d => n800, outb => 
                           n3334);
   U913 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_30_5_port, 
                           outb => n800);
   U914 : oai22 port map( a => n177, b => n796, c => n797, d => n801, outb => 
                           n3333);
   U915 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_30_4_port, 
                           outb => n801);
   U916 : oai22 port map( a => n175, b => n796, c => n797, d => n802, outb => 
                           n3332);
   U917 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_30_3_port, 
                           outb => n802);
   U918 : oai22 port map( a => n173, b => n796, c => n797, d => n803, outb => 
                           n3331);
   U919 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_30_2_port, 
                           outb => n803);
   U920 : oai22 port map( a => n171, b => n796, c => n797, d => n804, outb => 
                           n3330);
   U921 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_30_1_port, 
                           outb => n804);
   U922 : oai22 port map( a => n169, b => n796, c => n797, d => n805, outb => 
                           n3329);
   U923 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_30_0_port, 
                           outb => n805);
   U924 : oai22 port map( a => n183, b => n806, c => n807, d => n808, outb => 
                           n3328);
   U925 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_29_7_port, 
                           outb => n808);
   U926 : oai22 port map( a => n181, b => n806, c => n807, d => n809, outb => 
                           n3327);
   U927 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_29_6_port, 
                           outb => n809);
   U928 : oai22 port map( a => n179, b => n806, c => n807, d => n810, outb => 
                           n3326);
   U929 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_29_5_port, 
                           outb => n810);
   U930 : oai22 port map( a => n177, b => n806, c => n807, d => n811, outb => 
                           n3325);
   U931 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_29_4_port, 
                           outb => n811);
   U932 : oai22 port map( a => n175, b => n806, c => n807, d => n812, outb => 
                           n3324);
   U933 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_29_3_port, 
                           outb => n812);
   U934 : oai22 port map( a => n173, b => n806, c => n807, d => n813, outb => 
                           n3323);
   U935 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_29_2_port, 
                           outb => n813);
   U936 : oai22 port map( a => n171, b => n806, c => n807, d => n814, outb => 
                           n3322);
   U937 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_29_1_port, 
                           outb => n814);
   U938 : oai22 port map( a => n169, b => n806, c => n807, d => n815, outb => 
                           n3321);
   U939 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_29_0_port, 
                           outb => n815);
   U940 : oai22 port map( a => n183, b => n816, c => n817, d => n818, outb => 
                           n3320);
   U941 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_28_7_port, 
                           outb => n818);
   U942 : oai22 port map( a => n181, b => n816, c => n817, d => n819, outb => 
                           n3319);
   U943 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_28_6_port, 
                           outb => n819);
   U944 : oai22 port map( a => n179, b => n816, c => n817, d => n820, outb => 
                           n3318);
   U945 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_28_5_port, 
                           outb => n820);
   U946 : oai22 port map( a => n177, b => n816, c => n817, d => n821, outb => 
                           n3317);
   U947 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_28_4_port, 
                           outb => n821);
   U948 : oai22 port map( a => n175, b => n816, c => n817, d => n822, outb => 
                           n3316);
   U949 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_28_3_port, 
                           outb => n822);
   U950 : oai22 port map( a => n173, b => n816, c => n817, d => n823, outb => 
                           n3315);
   U951 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_28_2_port, 
                           outb => n823);
   U952 : oai22 port map( a => n171, b => n816, c => n817, d => n824, outb => 
                           n3314);
   U953 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_28_1_port, 
                           outb => n824);
   U954 : oai22 port map( a => n169, b => n816, c => n817, d => n825, outb => 
                           n3313);
   U955 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_28_0_port, 
                           outb => n825);
   U956 : oai22 port map( a => n183, b => n826, c => n827, d => n828, outb => 
                           n3312);
   U957 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_27_7_port, 
                           outb => n828);
   U958 : oai22 port map( a => n181, b => n826, c => n827, d => n829, outb => 
                           n3311);
   U959 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_27_6_port, 
                           outb => n829);
   U960 : oai22 port map( a => n179, b => n826, c => n827, d => n830, outb => 
                           n3310);
   U961 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_27_5_port, 
                           outb => n830);
   U962 : oai22 port map( a => n177, b => n826, c => n827, d => n831, outb => 
                           n3309);
   U963 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_27_4_port, 
                           outb => n831);
   U964 : oai22 port map( a => n175, b => n826, c => n827, d => n832, outb => 
                           n3308);
   U965 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_27_3_port, 
                           outb => n832);
   U966 : oai22 port map( a => n173, b => n826, c => n827, d => n833, outb => 
                           n3307);
   U967 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_27_2_port, 
                           outb => n833);
   U968 : oai22 port map( a => n171, b => n826, c => n827, d => n834, outb => 
                           n3306);
   U969 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_27_1_port, 
                           outb => n834);
   U970 : oai22 port map( a => n169, b => n826, c => n827, d => n835, outb => 
                           n3305);
   U971 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_27_0_port, 
                           outb => n835);
   U972 : oai22 port map( a => n183, b => n836, c => n837, d => n838, outb => 
                           n3304);
   U973 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_26_7_port, 
                           outb => n838);
   U974 : oai22 port map( a => n181, b => n836, c => n837, d => n839, outb => 
                           n3303);
   U975 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_26_6_port, 
                           outb => n839);
   U976 : oai22 port map( a => n179, b => n836, c => n837, d => n840, outb => 
                           n3302);
   U977 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_26_5_port, 
                           outb => n840);
   U978 : oai22 port map( a => n177, b => n836, c => n837, d => n841, outb => 
                           n3301);
   U979 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_26_4_port, 
                           outb => n841);
   U980 : oai22 port map( a => n175, b => n836, c => n837, d => n842, outb => 
                           n3300);
   U981 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_26_3_port, 
                           outb => n842);
   U982 : oai22 port map( a => n173, b => n836, c => n837, d => n843, outb => 
                           n3299);
   U983 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_26_2_port, 
                           outb => n843);
   U984 : oai22 port map( a => n171, b => n836, c => n837, d => n844, outb => 
                           n3298);
   U985 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_26_1_port, 
                           outb => n844);
   U986 : oai22 port map( a => n169, b => n836, c => n837, d => n845, outb => 
                           n3297);
   U987 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_26_0_port, 
                           outb => n845);
   U988 : oai22 port map( a => n183, b => n846, c => n847, d => n848, outb => 
                           n3296);
   U989 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_25_7_port, 
                           outb => n848);
   U990 : oai22 port map( a => n181, b => n846, c => n847, d => n849, outb => 
                           n3295);
   U991 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_25_6_port, 
                           outb => n849);
   U992 : oai22 port map( a => n179, b => n846, c => n847, d => n850, outb => 
                           n3294);
   U993 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_25_5_port, 
                           outb => n850);
   U994 : oai22 port map( a => n177, b => n846, c => n847, d => n851, outb => 
                           n3293);
   U995 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_25_4_port, 
                           outb => n851);
   U996 : oai22 port map( a => n175, b => n846, c => n847, d => n852, outb => 
                           n3292);
   U997 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_25_3_port, 
                           outb => n852);
   U998 : oai22 port map( a => n173, b => n846, c => n847, d => n853, outb => 
                           n3291);
   U999 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_25_2_port, 
                           outb => n853);
   U1000 : oai22 port map( a => n171, b => n846, c => n847, d => n854, outb => 
                           n3290);
   U1001 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_25_1_port,
                           outb => n854);
   U1002 : oai22 port map( a => n169, b => n846, c => n847, d => n855, outb => 
                           n3289);
   U1003 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_25_0_port,
                           outb => n855);
   U1004 : oai22 port map( a => n183, b => n856, c => n857, d => n858, outb => 
                           n3288);
   U1005 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_24_7_port,
                           outb => n858);
   U1006 : oai22 port map( a => n181, b => n856, c => n857, d => n859, outb => 
                           n3287);
   U1007 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_24_6_port,
                           outb => n859);
   U1008 : oai22 port map( a => n179, b => n856, c => n857, d => n860, outb => 
                           n3286);
   U1009 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_24_5_port,
                           outb => n860);
   U1010 : oai22 port map( a => n177, b => n856, c => n857, d => n861, outb => 
                           n3285);
   U1011 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_24_4_port,
                           outb => n861);
   U1012 : oai22 port map( a => n175, b => n856, c => n857, d => n862, outb => 
                           n3284);
   U1013 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_24_3_port,
                           outb => n862);
   U1014 : oai22 port map( a => n173, b => n856, c => n857, d => n863, outb => 
                           n3283);
   U1015 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_24_2_port,
                           outb => n863);
   U1016 : oai22 port map( a => n171, b => n856, c => n857, d => n864, outb => 
                           n3282);
   U1017 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_24_1_port,
                           outb => n864);
   U1018 : oai22 port map( a => n169, b => n856, c => n857, d => n865, outb => 
                           n3281);
   U1019 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_24_0_port,
                           outb => n865);
   U1020 : oai22 port map( a => n183, b => n866, c => n867, d => n868, outb => 
                           n3280);
   U1021 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_23_7_port,
                           outb => n868);
   U1022 : oai22 port map( a => n181, b => n866, c => n867, d => n869, outb => 
                           n3279);
   U1023 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_23_6_port,
                           outb => n869);
   U1024 : oai22 port map( a => n179, b => n866, c => n867, d => n870, outb => 
                           n3278);
   U1025 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_23_5_port,
                           outb => n870);
   U1026 : oai22 port map( a => n177, b => n866, c => n867, d => n871, outb => 
                           n3277);
   U1027 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_23_4_port,
                           outb => n871);
   U1028 : oai22 port map( a => n175, b => n866, c => n867, d => n872, outb => 
                           n3276);
   U1029 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_23_3_port,
                           outb => n872);
   U1030 : oai22 port map( a => n173, b => n866, c => n867, d => n873, outb => 
                           n3275);
   U1031 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_23_2_port,
                           outb => n873);
   U1032 : oai22 port map( a => n171, b => n866, c => n867, d => n874, outb => 
                           n3274);
   U1033 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_23_1_port,
                           outb => n874);
   U1034 : oai22 port map( a => n169, b => n866, c => n867, d => n875, outb => 
                           n3273);
   U1035 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_23_0_port,
                           outb => n875);
   U1036 : oai22 port map( a => n183, b => n876, c => n877, d => n878, outb => 
                           n3272);
   U1037 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_22_7_port,
                           outb => n878);
   U1038 : oai22 port map( a => n181, b => n876, c => n877, d => n879, outb => 
                           n3271);
   U1039 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_22_6_port,
                           outb => n879);
   U1040 : oai22 port map( a => n179, b => n876, c => n877, d => n880, outb => 
                           n3270);
   U1041 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_22_5_port,
                           outb => n880);
   U1042 : oai22 port map( a => n177, b => n876, c => n877, d => n881, outb => 
                           n3269);
   U1043 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_22_4_port,
                           outb => n881);
   U1044 : oai22 port map( a => n175, b => n876, c => n877, d => n882, outb => 
                           n3268);
   U1045 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_22_3_port,
                           outb => n882);
   U1046 : oai22 port map( a => n173, b => n876, c => n877, d => n883, outb => 
                           n3267);
   U1047 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_22_2_port,
                           outb => n883);
   U1048 : oai22 port map( a => n171, b => n876, c => n877, d => n884, outb => 
                           n3266);
   U1049 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_22_1_port,
                           outb => n884);
   U1050 : oai22 port map( a => n169, b => n876, c => n877, d => n885, outb => 
                           n3265);
   U1051 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_22_0_port,
                           outb => n885);
   U1052 : oai22 port map( a => n183, b => n886, c => n887, d => n524, outb => 
                           n3264);
   U1053 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_21_7_port,
                           outb => n524);
   U1054 : oai22 port map( a => n181, b => n886, c => n887, d => n563, outb => 
                           n3263);
   U1055 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_21_6_port,
                           outb => n563);
   U1056 : oai22 port map( a => n179, b => n886, c => n887, d => n598, outb => 
                           n3262);
   U1057 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_21_5_port,
                           outb => n598);
   U1058 : oai22 port map( a => n177, b => n886, c => n887, d => n633, outb => 
                           n3261);
   U1059 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_21_4_port,
                           outb => n633);
   U1060 : oai22 port map( a => n175, b => n886, c => n887, d => n667, outb => 
                           n3260);
   U1061 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_21_3_port,
                           outb => n667);
   U1062 : oai22 port map( a => n173, b => n886, c => n887, d => n701, outb => 
                           n3259);
   U1063 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_21_2_port,
                           outb => n701);
   U1064 : oai22 port map( a => n171, b => n886, c => n887, d => n735, outb => 
                           n3258);
   U1065 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_21_1_port,
                           outb => n735);
   U1066 : oai22 port map( a => n169, b => n886, c => n887, d => n769, outb => 
                           n3257);
   U1067 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_21_0_port,
                           outb => n769);
   U1068 : oai22 port map( a => n183, b => n888, c => n889, d => n526, outb => 
                           n3256);
   U1069 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_20_7_port,
                           outb => n526);
   U1070 : oai22 port map( a => n181, b => n888, c => n889, d => n564, outb => 
                           n3255);
   U1071 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_20_6_port,
                           outb => n564);
   U1072 : oai22 port map( a => n179, b => n888, c => n889, d => n599, outb => 
                           n3254);
   U1073 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_20_5_port,
                           outb => n599);
   U1074 : oai22 port map( a => n177, b => n888, c => n889, d => n634, outb => 
                           n3253);
   U1075 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_20_4_port,
                           outb => n634);
   U1076 : oai22 port map( a => n175, b => n888, c => n889, d => n668, outb => 
                           n3252);
   U1077 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_20_3_port,
                           outb => n668);
   U1078 : oai22 port map( a => n173, b => n888, c => n889, d => n702, outb => 
                           n3251);
   U1079 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_20_2_port,
                           outb => n702);
   U1080 : oai22 port map( a => n171, b => n888, c => n889, d => n736, outb => 
                           n3250);
   U1081 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_20_1_port,
                           outb => n736);
   U1082 : oai22 port map( a => n169, b => n888, c => n889, d => n770, outb => 
                           n3249);
   U1083 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_20_0_port,
                           outb => n770);
   U1084 : oai22 port map( a => n183, b => n890, c => n891, d => n528, outb => 
                           n3248);
   U1085 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_19_7_port,
                           outb => n528);
   U1086 : oai22 port map( a => n181, b => n890, c => n891, d => n565, outb => 
                           n3247);
   U1087 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_19_6_port,
                           outb => n565);
   U1088 : oai22 port map( a => n179, b => n890, c => n891, d => n600, outb => 
                           n3246);
   U1089 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_19_5_port,
                           outb => n600);
   U1090 : oai22 port map( a => n177, b => n890, c => n891, d => n635, outb => 
                           n3245);
   U1091 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_19_4_port,
                           outb => n635);
   U1092 : oai22 port map( a => n175, b => n890, c => n891, d => n669, outb => 
                           n3244);
   U1093 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_19_3_port,
                           outb => n669);
   U1094 : oai22 port map( a => n173, b => n890, c => n891, d => n703, outb => 
                           n3243);
   U1095 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_19_2_port,
                           outb => n703);
   U1096 : oai22 port map( a => n171, b => n890, c => n891, d => n737, outb => 
                           n3242);
   U1097 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_19_1_port,
                           outb => n737);
   U1098 : oai22 port map( a => n169, b => n890, c => n891, d => n771, outb => 
                           n3241);
   U1099 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_19_0_port,
                           outb => n771);
   U1100 : oai22 port map( a => n183, b => n892, c => n893, d => n894, outb => 
                           n3240);
   U1101 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_18_7_port,
                           outb => n894);
   U1102 : oai22 port map( a => n181, b => n892, c => n893, d => n895, outb => 
                           n3239);
   U1103 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_18_6_port,
                           outb => n895);
   U1104 : oai22 port map( a => n179, b => n892, c => n893, d => n896, outb => 
                           n3238);
   U1105 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_18_5_port,
                           outb => n896);
   U1106 : oai22 port map( a => n177, b => n892, c => n893, d => n897, outb => 
                           n3237);
   U1107 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_18_4_port,
                           outb => n897);
   U1108 : oai22 port map( a => n175, b => n892, c => n893, d => n898, outb => 
                           n3236);
   U1109 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_18_3_port,
                           outb => n898);
   U1110 : oai22 port map( a => n173, b => n892, c => n893, d => n899, outb => 
                           n3235);
   U1111 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_18_2_port,
                           outb => n899);
   U1112 : oai22 port map( a => n171, b => n892, c => n893, d => n900, outb => 
                           n3234);
   U1113 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_18_1_port,
                           outb => n900);
   U1114 : oai22 port map( a => n169, b => n892, c => n893, d => n901, outb => 
                           n3233);
   U1115 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_18_0_port,
                           outb => n901);
   U1116 : oai22 port map( a => n183, b => n902, c => n903, d => n904, outb => 
                           n3232);
   U1117 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_17_7_port,
                           outb => n904);
   U1118 : oai22 port map( a => n181, b => n902, c => n903, d => n905, outb => 
                           n3231);
   U1119 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_17_6_port,
                           outb => n905);
   U1120 : oai22 port map( a => n179, b => n902, c => n903, d => n906, outb => 
                           n3230);
   U1121 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_17_5_port,
                           outb => n906);
   U1122 : oai22 port map( a => n177, b => n902, c => n903, d => n907, outb => 
                           n3229);
   U1123 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_17_4_port,
                           outb => n907);
   U1124 : oai22 port map( a => n175, b => n902, c => n903, d => n908, outb => 
                           n3228);
   U1125 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_17_3_port,
                           outb => n908);
   U1126 : oai22 port map( a => n173, b => n902, c => n903, d => n909, outb => 
                           n3227);
   U1127 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_17_2_port,
                           outb => n909);
   U1128 : oai22 port map( a => n171, b => n902, c => n903, d => n910, outb => 
                           n3226);
   U1129 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_17_1_port,
                           outb => n910);
   U1130 : oai22 port map( a => n169, b => n902, c => n903, d => n911, outb => 
                           n3225);
   U1131 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_17_0_port,
                           outb => n911);
   U1132 : oai22 port map( a => n183, b => n912, c => n913, d => n914, outb => 
                           n3224);
   U1133 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_16_7_port,
                           outb => n914);
   U1134 : oai22 port map( a => n181, b => n912, c => n913, d => n915, outb => 
                           n3223);
   U1135 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_16_6_port,
                           outb => n915);
   U1136 : oai22 port map( a => n179, b => n912, c => n913, d => n916, outb => 
                           n3222);
   U1137 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_16_5_port,
                           outb => n916);
   U1138 : oai22 port map( a => n177, b => n912, c => n913, d => n917, outb => 
                           n3221);
   U1139 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_16_4_port,
                           outb => n917);
   U1140 : oai22 port map( a => n175, b => n912, c => n913, d => n918, outb => 
                           n3220);
   U1141 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_16_3_port,
                           outb => n918);
   U1142 : oai22 port map( a => n173, b => n912, c => n913, d => n919, outb => 
                           n3219);
   U1143 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_16_2_port,
                           outb => n919);
   U1144 : oai22 port map( a => n171, b => n912, c => n913, d => n920, outb => 
                           n3218);
   U1145 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_16_1_port,
                           outb => n920);
   U1146 : oai22 port map( a => n169, b => n912, c => n913, d => n921, outb => 
                           n3217);
   U1147 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_16_0_port,
                           outb => n921);
   U1148 : oai22 port map( a => n183, b => n922, c => n923, d => n924, outb => 
                           n3216);
   U1149 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_15_7_port,
                           outb => n924);
   U1150 : oai22 port map( a => n181, b => n922, c => n923, d => n925, outb => 
                           n3215);
   U1151 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_15_6_port,
                           outb => n925);
   U1152 : oai22 port map( a => n179, b => n922, c => n923, d => n926, outb => 
                           n3214);
   U1153 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_15_5_port,
                           outb => n926);
   U1154 : oai22 port map( a => n177, b => n922, c => n923, d => n927, outb => 
                           n3213);
   U1155 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_15_4_port,
                           outb => n927);
   U1156 : oai22 port map( a => n175, b => n922, c => n923, d => n928, outb => 
                           n3212);
   U1157 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_15_3_port,
                           outb => n928);
   U1158 : oai22 port map( a => n173, b => n922, c => n923, d => n929, outb => 
                           n3211);
   U1159 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_15_2_port,
                           outb => n929);
   U1160 : oai22 port map( a => n171, b => n922, c => n923, d => n930, outb => 
                           n3210);
   U1161 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_15_1_port,
                           outb => n930);
   U1162 : oai22 port map( a => n169, b => n922, c => n923, d => n931, outb => 
                           n3209);
   U1163 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_15_0_port,
                           outb => n931);
   U1164 : oai22 port map( a => n183, b => n932, c => n933, d => n934, outb => 
                           n3208);
   U1165 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_14_7_port,
                           outb => n934);
   U1166 : oai22 port map( a => n181, b => n932, c => n933, d => n935, outb => 
                           n3207);
   U1167 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_14_6_port,
                           outb => n935);
   U1168 : oai22 port map( a => n179, b => n932, c => n933, d => n936, outb => 
                           n3206);
   U1169 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_14_5_port,
                           outb => n936);
   U1170 : oai22 port map( a => n177, b => n932, c => n933, d => n937, outb => 
                           n3205);
   U1171 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_14_4_port,
                           outb => n937);
   U1172 : oai22 port map( a => n175, b => n932, c => n933, d => n938, outb => 
                           n3204);
   U1173 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_14_3_port,
                           outb => n938);
   U1174 : oai22 port map( a => n173, b => n932, c => n933, d => n939, outb => 
                           n3203);
   U1175 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_14_2_port,
                           outb => n939);
   U1176 : oai22 port map( a => n171, b => n932, c => n933, d => n940, outb => 
                           n3202);
   U1177 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_14_1_port,
                           outb => n940);
   U1178 : oai22 port map( a => n169, b => n932, c => n933, d => n941, outb => 
                           n3201);
   U1179 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_14_0_port,
                           outb => n941);
   U1180 : oai22 port map( a => n183, b => n942, c => n943, d => n536, outb => 
                           n3200);
   U1181 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_13_7_port,
                           outb => n536);
   U1182 : oai22 port map( a => n181, b => n942, c => n943, d => n572, outb => 
                           n3199);
   U1183 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_13_6_port,
                           outb => n572);
   U1184 : oai22 port map( a => n179, b => n942, c => n943, d => n607, outb => 
                           n3198);
   U1185 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_13_5_port,
                           outb => n607);
   U1186 : oai22 port map( a => n177, b => n942, c => n943, d => n642, outb => 
                           n3197);
   U1187 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_13_4_port,
                           outb => n642);
   U1188 : oai22 port map( a => n175, b => n942, c => n943, d => n676, outb => 
                           n3196);
   U1189 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_13_3_port,
                           outb => n676);
   U1190 : oai22 port map( a => n173, b => n942, c => n943, d => n710, outb => 
                           n3195);
   U1191 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_13_2_port,
                           outb => n710);
   U1192 : oai22 port map( a => n171, b => n942, c => n943, d => n744, outb => 
                           n3194);
   U1193 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_13_1_port,
                           outb => n744);
   U1194 : oai22 port map( a => n169, b => n942, c => n943, d => n778, outb => 
                           n3193);
   U1195 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_13_0_port,
                           outb => n778);
   U1196 : oai22 port map( a => n183, b => n944, c => n945, d => n537, outb => 
                           n3192);
   U1197 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_12_7_port,
                           outb => n537);
   U1198 : oai22 port map( a => n181, b => n944, c => n945, d => n573, outb => 
                           n3191);
   U1199 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_12_6_port,
                           outb => n573);
   U1200 : oai22 port map( a => n179, b => n944, c => n945, d => n608, outb => 
                           n3190);
   U1201 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_12_5_port,
                           outb => n608);
   U1202 : oai22 port map( a => n177, b => n944, c => n945, d => n643, outb => 
                           n3189);
   U1203 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_12_4_port,
                           outb => n643);
   U1204 : inv port map( inb => load_n_store_lazy_in_2_4_port, outb => n177);
   U1205 : oai22 port map( a => n175, b => n944, c => n945, d => n677, outb => 
                           n3188);
   U1206 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_12_3_port,
                           outb => n677);
   U1207 : inv port map( inb => load_n_store_lazy_in_2_3_port, outb => n175);
   U1208 : oai22 port map( a => n173, b => n944, c => n945, d => n711, outb => 
                           n3187);
   U1209 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_12_2_port,
                           outb => n711);
   U1210 : inv port map( inb => load_n_store_lazy_in_2_2_port, outb => n173);
   U1211 : oai22 port map( a => n171, b => n944, c => n945, d => n745, outb => 
                           n3186);
   U1212 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_12_1_port,
                           outb => n745);
   U1213 : inv port map( inb => load_n_store_lazy_in_2_1_port, outb => n171);
   U1214 : oai22 port map( a => n169, b => n944, c => n945, d => n779, outb => 
                           n3185);
   U1215 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_12_0_port,
                           outb => n779);
   U1216 : inv port map( inb => load_n_store_lazy_in_2_0_port, outb => n169);
   U1217 : oai22 port map( a => n183, b => n380, c => n381, d => n538, outb => 
                           n3184);
   U1218 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_11_7_port,
                           outb => n538);
   U1219 : inv port map( inb => load_n_store_lazy_in_2_7_port, outb => n183);
   U1220 : oai22 port map( a => n181, b => n380, c => n381, d => n574, outb => 
                           n3183);
   U1221 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_11_6_port,
                           outb => n574);
   U1222 : inv port map( inb => load_n_store_lazy_in_2_6_port, outb => n181);
   U1223 : oai22 port map( a => n179, b => n380, c => n381, d => n609, outb => 
                           n3182);
   U1224 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_11_5_port,
                           outb => n609);
   U1225 : inv port map( inb => load_n_store_lazy_in_2_5_port, outb => n179);
   U1226 : oai22 port map( a => n193, b => n380, c => n381, d => n946, outb => 
                           n2653);
   U1227 : oai22 port map( a => n191, b => n380, c => n381, d => n947, outb => 
                           n2652);
   U1228 : oai22 port map( a => n189, b => n380, c => n381, d => n948, outb => 
                           n2651);
   U1229 : oai22 port map( a => n187, b => n380, c => n381, d => n949, outb => 
                           n2650);
   U1230 : oai22 port map( a => n185, b => n380, c => n381, d => n950, outb => 
                           n2649);
   U1231 : oai22 port map( a => n199, b => n387, c => n388, d => n951, outb => 
                           n2648);
   U1232 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_10_7_port,
                           outb => n951);
   U1233 : oai22 port map( a => n197, b => n387, c => n388, d => n952, outb => 
                           n2647);
   U1234 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_10_6_port,
                           outb => n952);
   U1235 : oai22 port map( a => n195, b => n387, c => n388, d => n953, outb => 
                           n2646);
   U1236 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_10_5_port,
                           outb => n953);
   U1237 : oai22 port map( a => n193, b => n387, c => n388, d => n954, outb => 
                           n2645);
   U1238 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_10_4_port,
                           outb => n954);
   U1239 : oai22 port map( a => n191, b => n387, c => n388, d => n955, outb => 
                           n2644);
   U1240 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_10_3_port,
                           outb => n955);
   U1241 : oai22 port map( a => n189, b => n387, c => n388, d => n956, outb => 
                           n2643);
   U1242 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_10_2_port,
                           outb => n956);
   U1243 : oai22 port map( a => n187, b => n387, c => n388, d => n957, outb => 
                           n2642);
   U1244 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_10_1_port,
                           outb => n957);
   U1245 : oai22 port map( a => n185, b => n387, c => n388, d => n958, outb => 
                           n2641);
   U1246 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_10_0_port,
                           outb => n958);
   U1247 : oai22 port map( a => n199, b => n397, c => n398, d => n959, outb => 
                           n2640);
   U1248 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_9_7_port, 
                           outb => n959);
   U1249 : oai22 port map( a => n197, b => n397, c => n398, d => n960, outb => 
                           n2639);
   U1250 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_9_6_port, 
                           outb => n960);
   U1251 : oai22 port map( a => n195, b => n397, c => n398, d => n961, outb => 
                           n2638);
   U1252 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_9_5_port, 
                           outb => n961);
   U1253 : oai22 port map( a => n193, b => n397, c => n398, d => n962, outb => 
                           n2637);
   U1254 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_9_4_port, 
                           outb => n962);
   U1255 : oai22 port map( a => n191, b => n397, c => n398, d => n963, outb => 
                           n2636);
   U1256 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_9_3_port, 
                           outb => n963);
   U1257 : oai22 port map( a => n189, b => n397, c => n398, d => n964, outb => 
                           n2635);
   U1258 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_9_2_port, 
                           outb => n964);
   U1259 : oai22 port map( a => n187, b => n397, c => n398, d => n965, outb => 
                           n2634);
   U1260 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_9_1_port, 
                           outb => n965);
   U1261 : oai22 port map( a => n185, b => n397, c => n398, d => n966, outb => 
                           n2633);
   U1262 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_9_0_port, 
                           outb => n966);
   U1263 : oai22 port map( a => n199, b => n407, c => n408, d => n967, outb => 
                           n2632);
   U1264 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_8_7_port, 
                           outb => n967);
   U1265 : oai22 port map( a => n197, b => n407, c => n408, d => n968, outb => 
                           n2631);
   U1266 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_8_6_port, 
                           outb => n968);
   U1267 : oai22 port map( a => n195, b => n407, c => n408, d => n969, outb => 
                           n2630);
   U1268 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_8_5_port, 
                           outb => n969);
   U1269 : oai22 port map( a => n193, b => n407, c => n408, d => n970, outb => 
                           n2629);
   U1270 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_8_4_port, 
                           outb => n970);
   U1271 : oai22 port map( a => n191, b => n407, c => n408, d => n971, outb => 
                           n2628);
   U1272 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_8_3_port, 
                           outb => n971);
   U1273 : oai22 port map( a => n189, b => n407, c => n408, d => n972, outb => 
                           n2627);
   U1274 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_8_2_port, 
                           outb => n972);
   U1275 : oai22 port map( a => n187, b => n407, c => n408, d => n973, outb => 
                           n2626);
   U1276 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_8_1_port, 
                           outb => n973);
   U1277 : oai22 port map( a => n185, b => n407, c => n408, d => n974, outb => 
                           n2625);
   U1278 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_8_0_port, 
                           outb => n974);
   U1279 : oai22 port map( a => n199, b => n417, c => n418, d => n975, outb => 
                           n2624);
   U1280 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_7_7_port, 
                           outb => n975);
   U1281 : oai22 port map( a => n197, b => n417, c => n418, d => n976, outb => 
                           n2623);
   U1282 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_7_6_port, 
                           outb => n976);
   U1283 : oai22 port map( a => n195, b => n417, c => n418, d => n977, outb => 
                           n2622);
   U1284 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_7_5_port, 
                           outb => n977);
   U1285 : oai22 port map( a => n193, b => n417, c => n418, d => n978, outb => 
                           n2621);
   U1286 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_7_4_port, 
                           outb => n978);
   U1287 : oai22 port map( a => n191, b => n417, c => n418, d => n979, outb => 
                           n2620);
   U1288 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_7_3_port, 
                           outb => n979);
   U1289 : oai22 port map( a => n189, b => n417, c => n418, d => n980, outb => 
                           n2619);
   U1290 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_7_2_port, 
                           outb => n980);
   U1291 : oai22 port map( a => n187, b => n417, c => n418, d => n981, outb => 
                           n2618);
   U1292 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_7_1_port, 
                           outb => n981);
   U1293 : oai22 port map( a => n185, b => n417, c => n418, d => n982, outb => 
                           n2617);
   U1294 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_7_0_port, 
                           outb => n982);
   U1295 : oai22 port map( a => n199, b => n427, c => n428, d => n983, outb => 
                           n2616);
   U1296 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_6_7_port, 
                           outb => n983);
   U1297 : oai22 port map( a => n197, b => n427, c => n428, d => n984, outb => 
                           n2615);
   U1298 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_6_6_port, 
                           outb => n984);
   U1299 : oai22 port map( a => n195, b => n427, c => n428, d => n985, outb => 
                           n2614);
   U1300 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_6_5_port, 
                           outb => n985);
   U1301 : oai22 port map( a => n193, b => n427, c => n428, d => n986, outb => 
                           n2613);
   U1302 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_6_4_port, 
                           outb => n986);
   U1303 : oai22 port map( a => n191, b => n427, c => n428, d => n987, outb => 
                           n2612);
   U1304 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_6_3_port, 
                           outb => n987);
   U1305 : oai22 port map( a => n189, b => n427, c => n428, d => n988, outb => 
                           n2611);
   U1306 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_6_2_port, 
                           outb => n988);
   U1307 : oai22 port map( a => n187, b => n427, c => n428, d => n989, outb => 
                           n2610);
   U1308 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_6_1_port, 
                           outb => n989);
   U1309 : oai22 port map( a => n185, b => n427, c => n428, d => n990, outb => 
                           n2609);
   U1310 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_6_0_port, 
                           outb => n990);
   U1311 : oai22 port map( a => n199, b => n437, c => n438, d => n991, outb => 
                           n2608);
   U1312 : oai22 port map( a => n197, b => n437, c => n438, d => n992, outb => 
                           n2607);
   U1313 : oai22 port map( a => n195, b => n437, c => n438, d => n993, outb => 
                           n2606);
   U1314 : oai22 port map( a => n193, b => n437, c => n438, d => n994, outb => 
                           n2605);
   U1315 : oai22 port map( a => n191, b => n437, c => n438, d => n995, outb => 
                           n2604);
   U1316 : oai22 port map( a => n189, b => n437, c => n438, d => n996, outb => 
                           n2603);
   U1317 : oai22 port map( a => n187, b => n437, c => n438, d => n997, outb => 
                           n2602);
   U1318 : oai22 port map( a => n185, b => n437, c => n438, d => n998, outb => 
                           n2601);
   U1319 : oai22 port map( a => n199, b => n447, c => n448, d => n999, outb => 
                           n2600);
   U1320 : oai22 port map( a => n197, b => n447, c => n448, d => n1000, outb =>
                           n2599);
   U1321 : oai22 port map( a => n195, b => n447, c => n448, d => n1001, outb =>
                           n2598);
   U1322 : oai22 port map( a => n193, b => n447, c => n448, d => n1002, outb =>
                           n2597);
   U1323 : oai22 port map( a => n191, b => n447, c => n448, d => n1003, outb =>
                           n2596);
   U1324 : oai22 port map( a => n189, b => n447, c => n448, d => n1004, outb =>
                           n2595);
   U1325 : oai22 port map( a => n187, b => n447, c => n448, d => n1005, outb =>
                           n2594);
   U1326 : oai22 port map( a => n185, b => n447, c => n448, d => n1006, outb =>
                           n2593);
   U1327 : oai22 port map( a => n199, b => n457, c => n458, d => n1007, outb =>
                           n2592);
   U1328 : oai22 port map( a => n197, b => n457, c => n458, d => n1008, outb =>
                           n2591);
   U1329 : oai22 port map( a => n195, b => n457, c => n458, d => n1009, outb =>
                           n2590);
   U1330 : oai22 port map( a => n193, b => n457, c => n458, d => n1010, outb =>
                           n2589);
   U1331 : oai22 port map( a => n191, b => n457, c => n458, d => n1011, outb =>
                           n2588);
   U1332 : oai22 port map( a => n189, b => n457, c => n458, d => n1012, outb =>
                           n2587);
   U1333 : oai22 port map( a => n187, b => n457, c => n458, d => n1013, outb =>
                           n2586);
   U1334 : oai22 port map( a => n185, b => n457, c => n458, d => n1014, outb =>
                           n2585);
   U1335 : oai22 port map( a => n199, b => n467, c => n468, d => n1015, outb =>
                           n2584);
   U1336 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_2_7_port, 
                           outb => n1015);
   U1337 : oai22 port map( a => n197, b => n467, c => n468, d => n1016, outb =>
                           n2583);
   U1338 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_2_6_port, 
                           outb => n1016);
   U1339 : oai22 port map( a => n195, b => n467, c => n468, d => n1017, outb =>
                           n2582);
   U1340 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_2_5_port, 
                           outb => n1017);
   U1341 : oai22 port map( a => n193, b => n467, c => n468, d => n1018, outb =>
                           n2581);
   U1342 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_2_4_port, 
                           outb => n1018);
   U1343 : oai22 port map( a => n191, b => n467, c => n468, d => n1019, outb =>
                           n2580);
   U1344 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_2_3_port, 
                           outb => n1019);
   U1345 : oai22 port map( a => n189, b => n467, c => n468, d => n1020, outb =>
                           n2579);
   U1346 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_2_2_port, 
                           outb => n1020);
   U1347 : oai22 port map( a => n187, b => n467, c => n468, d => n1021, outb =>
                           n2578);
   U1348 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_2_1_port, 
                           outb => n1021);
   U1349 : oai22 port map( a => n185, b => n467, c => n468, d => n1022, outb =>
                           n2577);
   U1350 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_2_0_port, 
                           outb => n1022);
   U1351 : oai22 port map( a => n199, b => n477, c => n478, d => n1023, outb =>
                           n2576);
   U1352 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_1_7_port, 
                           outb => n1023);
   U1353 : oai22 port map( a => n197, b => n477, c => n478, d => n1024, outb =>
                           n2575);
   U1354 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_1_6_port, 
                           outb => n1024);
   U1355 : oai22 port map( a => n195, b => n477, c => n478, d => n1025, outb =>
                           n2574);
   U1356 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_1_5_port, 
                           outb => n1025);
   U1357 : oai22 port map( a => n193, b => n477, c => n478, d => n1026, outb =>
                           n2573);
   U1358 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_1_4_port, 
                           outb => n1026);
   U1359 : oai22 port map( a => n191, b => n477, c => n478, d => n1027, outb =>
                           n2572);
   U1360 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_1_3_port, 
                           outb => n1027);
   U1361 : oai22 port map( a => n189, b => n477, c => n478, d => n1028, outb =>
                           n2571);
   U1362 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_1_2_port, 
                           outb => n1028);
   U1363 : oai22 port map( a => n187, b => n477, c => n478, d => n1029, outb =>
                           n2570);
   U1364 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_1_1_port, 
                           outb => n1029);
   U1365 : oai22 port map( a => n185, b => n477, c => n478, d => n1030, outb =>
                           n2569);
   U1366 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_1_0_port, 
                           outb => n1030);
   U1367 : oai22 port map( a => n199, b => n487, c => n488, d => n1031, outb =>
                           n2568);
   U1368 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_0_7_port, 
                           outb => n1031);
   U1369 : oai22 port map( a => n197, b => n487, c => n488, d => n1032, outb =>
                           n2567);
   U1370 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_0_6_port, 
                           outb => n1032);
   U1371 : oai22 port map( a => n195, b => n487, c => n488, d => n1033, outb =>
                           n2566);
   U1372 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_0_5_port, 
                           outb => n1033);
   U1373 : oai22 port map( a => n193, b => n487, c => n488, d => n1034, outb =>
                           n2565);
   U1374 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_0_4_port, 
                           outb => n1034);
   U1375 : oai22 port map( a => n191, b => n487, c => n488, d => n1035, outb =>
                           n2564);
   U1376 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_0_3_port, 
                           outb => n1035);
   U1377 : oai22 port map( a => n189, b => n487, c => n488, d => n1036, outb =>
                           n2563);
   U1378 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_0_2_port, 
                           outb => n1036);
   U1379 : oai22 port map( a => n187, b => n487, c => n488, d => n1037, outb =>
                           n2562);
   U1380 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_0_1_port, 
                           outb => n1037);
   U1381 : oai22 port map( a => n185, b => n487, c => n488, d => n1038, outb =>
                           n2561);
   U1382 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_0_0_port, 
                           outb => n1038);
   U1383 : nand4 port map( a => n1039, b => n1040, c => n1041, d => n1042, outb
                           => n2311);
   U1384 : aoi22 port map( a => n1043, b => n1044, c => load_n_store_we_i, d =>
                           load_n_store_lazy_in_1_7_port, outb => n1042);
   U1385 : nor3 port map( a => n1045, b => n1046, c => n1047, outb => n1044);
   U1386 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_26_7_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_31_7_port, d =>
                           n370, outb => n1047);
   U1387 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_25_7_port, 
                           b => n507, outb => n1046);
   U1388 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_30_7_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_24_7_port, d =>
                           n509, outb => n1045);
   U1389 : nor3 port map( a => n1048, b => n1049, c => n512, outb => n1043);
   U1390 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_27_7_port, 
                           b => n513, outb => n1049);
   U1391 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_28_7_port,
                           b => n514, c => 
                           load_n_store_RGB_Array_1_block_ram_r_29_7_port, d =>
                           n515, outb => n1048);
   U1392 : nand4 port map( a => n516, b => n1050, c => n1051, d => n1052, outb 
                           => n1041);
   U1393 : nor3 port map( a => n1053, b => n1054, c => n1055, outb => n1052);
   U1394 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_18_7_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_23_7_port, d =>
                           n370, outb => n1055);
   U1395 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_17_7_port, 
                           b => n507, outb => n1054);
   U1396 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_22_7_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_16_7_port, d =>
                           n509, outb => n1053);
   U1397 : aoi22 port map( a => n523, b => n1056, c => n525, d => n1057, outb 
                           => n1051);
   U1398 : nand2 port map( a => n527, b => n1058, outb => n1050);
   U1399 : nand4 port map( a => n529, b => n1059, c => n1060, d => n1061, outb 
                           => n1040);
   U1400 : nor3 port map( a => n1062, b => n1063, c => n1064, outb => n1061);
   U1401 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_10_7_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_15_7_port, d =>
                           n370, outb => n1064);
   U1402 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_9_7_port, b
                           => n507, outb => n1063);
   U1403 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_14_7_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_8_7_port, d => 
                           n509, outb => n1062);
   U1404 : aoi22 port map( a => n523, b => n1065, c => n525, d => n1066, outb 
                           => n1060);
   U1405 : nand2 port map( a => n527, b => n1067, outb => n1059);
   U1406 : nand4 port map( a => n539, b => n1068, c => n1069, d => n1070, outb 
                           => n1039);
   U1407 : nor3 port map( a => n1071, b => n1072, c => n1073, outb => n1070);
   U1408 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_2_7_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_7_7_port, d => 
                           n370, outb => n1073);
   U1409 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_1_7_port, b
                           => n507, outb => n1072);
   U1410 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_6_7_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_0_7_port, d => 
                           n509, outb => n1071);
   U1411 : aoi22 port map( a => n523, b => n991, c => n525, d => n999, outb => 
                           n1069);
   U1412 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_4_7_port, 
                           outb => n999);
   U1413 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_5_7_port, 
                           outb => n991);
   U1414 : nand2 port map( a => n527, b => n1007, outb => n1068);
   U1415 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_3_7_port, 
                           outb => n1007);
   U1416 : nand4 port map( a => n1074, b => n1075, c => n1076, d => n1077, outb
                           => n2308);
   U1417 : aoi22 port map( a => n1078, b => n1079, c => load_n_store_we_i, d =>
                           load_n_store_lazy_in_1_6_port, outb => n1077);
   U1418 : nor3 port map( a => n1080, b => n1081, c => n1082, outb => n1079);
   U1419 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_26_6_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_31_6_port, d =>
                           n370, outb => n1082);
   U1420 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_25_6_port, 
                           b => n507, outb => n1081);
   U1421 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_30_6_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_24_6_port, d =>
                           n509, outb => n1080);
   U1422 : nor3 port map( a => n1083, b => n1084, c => n512, outb => n1078);
   U1423 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_27_6_port, 
                           b => n513, outb => n1084);
   U1424 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_28_6_port,
                           b => n514, c => 
                           load_n_store_RGB_Array_1_block_ram_r_29_6_port, d =>
                           n515, outb => n1083);
   U1425 : nand4 port map( a => n516, b => n1085, c => n1086, d => n1087, outb 
                           => n1076);
   U1426 : nor3 port map( a => n1088, b => n1089, c => n1090, outb => n1087);
   U1427 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_18_6_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_23_6_port, d =>
                           n370, outb => n1090);
   U1428 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_17_6_port, 
                           b => n507, outb => n1089);
   U1429 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_22_6_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_16_6_port, d =>
                           n509, outb => n1088);
   U1430 : aoi22 port map( a => n523, b => n1091, c => n525, d => n1092, outb 
                           => n1086);
   U1431 : nand2 port map( a => n527, b => n1093, outb => n1085);
   U1432 : nand4 port map( a => n529, b => n1094, c => n1095, d => n1096, outb 
                           => n1075);
   U1433 : nor3 port map( a => n1097, b => n1098, c => n1099, outb => n1096);
   U1434 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_10_6_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_15_6_port, d =>
                           n370, outb => n1099);
   U1435 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_9_6_port, b
                           => n507, outb => n1098);
   U1436 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_14_6_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_8_6_port, d => 
                           n509, outb => n1097);
   U1437 : aoi22 port map( a => n523, b => n1100, c => n525, d => n1101, outb 
                           => n1095);
   U1438 : nand2 port map( a => n527, b => n1102, outb => n1094);
   U1439 : nand4 port map( a => n539, b => n1103, c => n1104, d => n1105, outb 
                           => n1074);
   U1440 : nor3 port map( a => n1106, b => n1107, c => n1108, outb => n1105);
   U1441 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_2_6_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_7_6_port, d => 
                           n370, outb => n1108);
   U1442 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_1_6_port, b
                           => n507, outb => n1107);
   U1443 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_6_6_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_0_6_port, d => 
                           n509, outb => n1106);
   U1444 : aoi22 port map( a => n523, b => n992, c => n525, d => n1000, outb =>
                           n1104);
   U1445 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_4_6_port, 
                           outb => n1000);
   U1446 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_5_6_port, 
                           outb => n992);
   U1447 : nand2 port map( a => n527, b => n1008, outb => n1103);
   U1448 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_3_6_port, 
                           outb => n1008);
   U1449 : nand4 port map( a => n1109, b => n1110, c => n1111, d => n1112, outb
                           => n2305);
   U1450 : aoi22 port map( a => n1113, b => n1114, c => load_n_store_we_i, d =>
                           load_n_store_lazy_in_1_5_port, outb => n1112);
   U1451 : nor3 port map( a => n1115, b => n1116, c => n1117, outb => n1114);
   U1452 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_26_5_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_31_5_port, d =>
                           n370, outb => n1117);
   U1453 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_25_5_port, 
                           b => n507, outb => n1116);
   U1454 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_30_5_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_24_5_port, d =>
                           n509, outb => n1115);
   U1455 : nor3 port map( a => n1118, b => n1119, c => n512, outb => n1113);
   U1456 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_27_5_port, 
                           b => n513, outb => n1119);
   U1457 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_28_5_port,
                           b => n514, c => 
                           load_n_store_RGB_Array_1_block_ram_r_29_5_port, d =>
                           n515, outb => n1118);
   U1458 : nand4 port map( a => n516, b => n1120, c => n1121, d => n1122, outb 
                           => n1111);
   U1459 : nor3 port map( a => n1123, b => n1124, c => n1125, outb => n1122);
   U1460 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_18_5_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_23_5_port, d =>
                           n370, outb => n1125);
   U1461 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_17_5_port, 
                           b => n507, outb => n1124);
   U1462 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_22_5_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_16_5_port, d =>
                           n509, outb => n1123);
   U1463 : aoi22 port map( a => n523, b => n1126, c => n525, d => n1127, outb 
                           => n1121);
   U1464 : nand2 port map( a => n527, b => n1128, outb => n1120);
   U1465 : nand4 port map( a => n529, b => n1129, c => n1130, d => n1131, outb 
                           => n1110);
   U1466 : nor3 port map( a => n1132, b => n1133, c => n1134, outb => n1131);
   U1467 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_10_5_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_15_5_port, d =>
                           n370, outb => n1134);
   U1468 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_9_5_port, b
                           => n507, outb => n1133);
   U1469 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_14_5_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_8_5_port, d => 
                           n509, outb => n1132);
   U1470 : aoi22 port map( a => n523, b => n1135, c => n525, d => n1136, outb 
                           => n1130);
   U1471 : nand2 port map( a => n527, b => n1137, outb => n1129);
   U1472 : nand4 port map( a => n539, b => n1138, c => n1139, d => n1140, outb 
                           => n1109);
   U1473 : nor3 port map( a => n1141, b => n1142, c => n1143, outb => n1140);
   U1474 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_2_5_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_7_5_port, d => 
                           n370, outb => n1143);
   U1475 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_1_5_port, b
                           => n507, outb => n1142);
   U1476 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_6_5_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_0_5_port, d => 
                           n509, outb => n1141);
   U1477 : aoi22 port map( a => n523, b => n993, c => n525, d => n1001, outb =>
                           n1139);
   U1478 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_4_5_port, 
                           outb => n1001);
   U1479 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_5_5_port, 
                           outb => n993);
   U1480 : nand2 port map( a => n527, b => n1009, outb => n1138);
   U1481 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_3_5_port, 
                           outb => n1009);
   U1482 : nand4 port map( a => n1144, b => n1145, c => n1146, d => n1147, outb
                           => n2302);
   U1483 : aoi22 port map( a => n1148, b => n1149, c => load_n_store_we_i, d =>
                           load_n_store_lazy_in_1_4_port, outb => n1147);
   U1484 : nor3 port map( a => n1150, b => n1151, c => n1152, outb => n1149);
   U1485 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_26_4_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_31_4_port, d =>
                           n370, outb => n1152);
   U1486 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_25_4_port, 
                           b => n507, outb => n1151);
   U1487 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_30_4_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_24_4_port, d =>
                           n509, outb => n1150);
   U1488 : nor3 port map( a => n1153, b => n1154, c => n512, outb => n1148);
   U1489 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_27_4_port, 
                           b => n513, outb => n1154);
   U1490 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_28_4_port,
                           b => n514, c => 
                           load_n_store_RGB_Array_1_block_ram_r_29_4_port, d =>
                           n515, outb => n1153);
   U1491 : nand4 port map( a => n516, b => n1155, c => n1156, d => n1157, outb 
                           => n1146);
   U1492 : nor3 port map( a => n1158, b => n1159, c => n1160, outb => n1157);
   U1493 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_18_4_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_23_4_port, d =>
                           n370, outb => n1160);
   U1494 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_17_4_port, 
                           b => n507, outb => n1159);
   U1495 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_22_4_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_16_4_port, d =>
                           n509, outb => n1158);
   U1496 : aoi22 port map( a => n523, b => n1161, c => n525, d => n1162, outb 
                           => n1156);
   U1497 : nand2 port map( a => n527, b => n1163, outb => n1155);
   U1498 : nand4 port map( a => n529, b => n1164, c => n1165, d => n1166, outb 
                           => n1145);
   U1499 : nor3 port map( a => n1167, b => n1168, c => n1169, outb => n1166);
   U1500 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_10_4_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_15_4_port, d =>
                           n370, outb => n1169);
   U1501 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_9_4_port, b
                           => n507, outb => n1168);
   U1502 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_14_4_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_8_4_port, d => 
                           n509, outb => n1167);
   U1503 : aoi22 port map( a => n523, b => n1170, c => n525, d => n1171, outb 
                           => n1165);
   U1504 : nand2 port map( a => n527, b => n946, outb => n1164);
   U1505 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_11_4_port,
                           outb => n946);
   U1506 : nand4 port map( a => n539, b => n1172, c => n1173, d => n1174, outb 
                           => n1144);
   U1507 : nor3 port map( a => n1175, b => n1176, c => n1177, outb => n1174);
   U1508 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_2_4_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_7_4_port, d => 
                           n370, outb => n1177);
   U1509 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_1_4_port, b
                           => n507, outb => n1176);
   U1510 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_6_4_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_0_4_port, d => 
                           n509, outb => n1175);
   U1511 : aoi22 port map( a => n523, b => n994, c => n525, d => n1002, outb =>
                           n1173);
   U1512 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_4_4_port, 
                           outb => n1002);
   U1513 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_5_4_port, 
                           outb => n994);
   U1514 : nand2 port map( a => n527, b => n1010, outb => n1172);
   U1515 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_3_4_port, 
                           outb => n1010);
   U1516 : nand4 port map( a => n1178, b => n1179, c => n1180, d => n1181, outb
                           => n2299);
   U1517 : aoi22 port map( a => n1182, b => n1183, c => load_n_store_we_i, d =>
                           load_n_store_lazy_in_1_3_port, outb => n1181);
   U1518 : nor3 port map( a => n1184, b => n1185, c => n1186, outb => n1183);
   U1519 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_26_3_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_31_3_port, d =>
                           n370, outb => n1186);
   U1520 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_25_3_port, 
                           b => n507, outb => n1185);
   U1521 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_30_3_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_24_3_port, d =>
                           n509, outb => n1184);
   U1522 : nor3 port map( a => n1187, b => n1188, c => n512, outb => n1182);
   U1523 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_27_3_port, 
                           b => n513, outb => n1188);
   U1524 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_28_3_port,
                           b => n514, c => 
                           load_n_store_RGB_Array_1_block_ram_r_29_3_port, d =>
                           n515, outb => n1187);
   U1525 : nand4 port map( a => n516, b => n1189, c => n1190, d => n1191, outb 
                           => n1180);
   U1526 : nor3 port map( a => n1192, b => n1193, c => n1194, outb => n1191);
   U1527 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_18_3_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_23_3_port, d =>
                           n370, outb => n1194);
   U1528 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_17_3_port, 
                           b => n507, outb => n1193);
   U1529 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_22_3_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_16_3_port, d =>
                           n509, outb => n1192);
   U1530 : aoi22 port map( a => n523, b => n1195, c => n525, d => n1196, outb 
                           => n1190);
   U1531 : nand2 port map( a => n527, b => n1197, outb => n1189);
   U1532 : nand4 port map( a => n529, b => n1198, c => n1199, d => n1200, outb 
                           => n1179);
   U1533 : nor3 port map( a => n1201, b => n1202, c => n1203, outb => n1200);
   U1534 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_10_3_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_15_3_port, d =>
                           n370, outb => n1203);
   U1535 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_9_3_port, b
                           => n507, outb => n1202);
   U1536 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_14_3_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_8_3_port, d => 
                           n509, outb => n1201);
   U1537 : aoi22 port map( a => n523, b => n1204, c => n525, d => n1205, outb 
                           => n1199);
   U1538 : nand2 port map( a => n527, b => n947, outb => n1198);
   U1539 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_11_3_port,
                           outb => n947);
   U1540 : nand4 port map( a => n539, b => n1206, c => n1207, d => n1208, outb 
                           => n1178);
   U1541 : nor3 port map( a => n1209, b => n1210, c => n1211, outb => n1208);
   U1542 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_2_3_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_7_3_port, d => 
                           n370, outb => n1211);
   U1543 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_1_3_port, b
                           => n507, outb => n1210);
   U1544 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_6_3_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_0_3_port, d => 
                           n509, outb => n1209);
   U1545 : aoi22 port map( a => n523, b => n995, c => n525, d => n1003, outb =>
                           n1207);
   U1546 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_4_3_port, 
                           outb => n1003);
   U1547 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_5_3_port, 
                           outb => n995);
   U1548 : nand2 port map( a => n527, b => n1011, outb => n1206);
   U1549 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_3_3_port, 
                           outb => n1011);
   U1550 : nand4 port map( a => n1212, b => n1213, c => n1214, d => n1215, outb
                           => n2296);
   U1551 : aoi22 port map( a => n1216, b => n1217, c => load_n_store_we_i, d =>
                           load_n_store_lazy_in_1_2_port, outb => n1215);
   U1552 : nor3 port map( a => n1218, b => n1219, c => n1220, outb => n1217);
   U1553 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_26_2_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_31_2_port, d =>
                           n370, outb => n1220);
   U1554 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_25_2_port, 
                           b => n507, outb => n1219);
   U1555 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_30_2_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_24_2_port, d =>
                           n509, outb => n1218);
   U1556 : nor3 port map( a => n1221, b => n1222, c => n512, outb => n1216);
   U1557 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_27_2_port, 
                           b => n513, outb => n1222);
   U1558 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_28_2_port,
                           b => n514, c => 
                           load_n_store_RGB_Array_1_block_ram_r_29_2_port, d =>
                           n515, outb => n1221);
   U1559 : nand4 port map( a => n516, b => n1223, c => n1224, d => n1225, outb 
                           => n1214);
   U1560 : nor3 port map( a => n1226, b => n1227, c => n1228, outb => n1225);
   U1561 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_18_2_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_23_2_port, d =>
                           n370, outb => n1228);
   U1562 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_17_2_port, 
                           b => n507, outb => n1227);
   U1563 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_22_2_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_16_2_port, d =>
                           n509, outb => n1226);
   U1564 : aoi22 port map( a => n523, b => n1229, c => n525, d => n1230, outb 
                           => n1224);
   U1565 : nand2 port map( a => n527, b => n1231, outb => n1223);
   U1566 : nand4 port map( a => n529, b => n1232, c => n1233, d => n1234, outb 
                           => n1213);
   U1567 : nor3 port map( a => n1235, b => n1236, c => n1237, outb => n1234);
   U1568 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_10_2_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_15_2_port, d =>
                           n370, outb => n1237);
   U1569 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_9_2_port, b
                           => n507, outb => n1236);
   U1570 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_14_2_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_8_2_port, d => 
                           n509, outb => n1235);
   U1571 : aoi22 port map( a => n523, b => n1238, c => n525, d => n1239, outb 
                           => n1233);
   U1572 : nand2 port map( a => n527, b => n948, outb => n1232);
   U1573 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_11_2_port,
                           outb => n948);
   U1574 : nand4 port map( a => n539, b => n1240, c => n1241, d => n1242, outb 
                           => n1212);
   U1575 : nor3 port map( a => n1243, b => n1244, c => n1245, outb => n1242);
   U1576 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_2_2_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_7_2_port, d => 
                           n370, outb => n1245);
   U1577 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_1_2_port, b
                           => n507, outb => n1244);
   U1578 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_6_2_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_0_2_port, d => 
                           n509, outb => n1243);
   U1579 : aoi22 port map( a => n523, b => n996, c => n525, d => n1004, outb =>
                           n1241);
   U1580 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_4_2_port, 
                           outb => n1004);
   U1581 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_5_2_port, 
                           outb => n996);
   U1582 : nand2 port map( a => n527, b => n1012, outb => n1240);
   U1583 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_3_2_port, 
                           outb => n1012);
   U1584 : nand4 port map( a => n1246, b => n1247, c => n1248, d => n1249, outb
                           => n2293);
   U1585 : aoi22 port map( a => n1250, b => n1251, c => load_n_store_we_i, d =>
                           load_n_store_lazy_in_1_1_port, outb => n1249);
   U1586 : nor3 port map( a => n1252, b => n1253, c => n1254, outb => n1251);
   U1587 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_26_1_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_31_1_port, d =>
                           n370, outb => n1254);
   U1588 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_25_1_port, 
                           b => n507, outb => n1253);
   U1589 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_30_1_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_24_1_port, d =>
                           n509, outb => n1252);
   U1590 : nor3 port map( a => n1255, b => n1256, c => n512, outb => n1250);
   U1591 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_27_1_port, 
                           b => n513, outb => n1256);
   U1592 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_28_1_port,
                           b => n514, c => 
                           load_n_store_RGB_Array_1_block_ram_r_29_1_port, d =>
                           n515, outb => n1255);
   U1593 : nand4 port map( a => n516, b => n1257, c => n1258, d => n1259, outb 
                           => n1248);
   U1594 : nor3 port map( a => n1260, b => n1261, c => n1262, outb => n1259);
   U1595 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_18_1_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_23_1_port, d =>
                           n370, outb => n1262);
   U1596 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_17_1_port, 
                           b => n507, outb => n1261);
   U1597 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_22_1_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_16_1_port, d =>
                           n509, outb => n1260);
   U1598 : aoi22 port map( a => n523, b => n1263, c => n525, d => n1264, outb 
                           => n1258);
   U1599 : nand2 port map( a => n527, b => n1265, outb => n1257);
   U1600 : nand4 port map( a => n529, b => n1266, c => n1267, d => n1268, outb 
                           => n1247);
   U1601 : nor3 port map( a => n1269, b => n1270, c => n1271, outb => n1268);
   U1602 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_10_1_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_15_1_port, d =>
                           n370, outb => n1271);
   U1603 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_9_1_port, b
                           => n507, outb => n1270);
   U1604 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_14_1_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_8_1_port, d => 
                           n509, outb => n1269);
   U1605 : aoi22 port map( a => n523, b => n1272, c => n525, d => n1273, outb 
                           => n1267);
   U1606 : nand2 port map( a => n527, b => n949, outb => n1266);
   U1607 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_11_1_port,
                           outb => n949);
   U1608 : nand4 port map( a => n539, b => n1274, c => n1275, d => n1276, outb 
                           => n1246);
   U1609 : nor3 port map( a => n1277, b => n1278, c => n1279, outb => n1276);
   U1610 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_2_1_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_7_1_port, d => 
                           n370, outb => n1279);
   U1611 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_1_1_port, b
                           => n507, outb => n1278);
   U1612 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_6_1_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_0_1_port, d => 
                           n509, outb => n1277);
   U1613 : aoi22 port map( a => n523, b => n997, c => n525, d => n1005, outb =>
                           n1275);
   U1614 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_4_1_port, 
                           outb => n1005);
   U1615 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_5_1_port, 
                           outb => n997);
   U1616 : nand2 port map( a => n527, b => n1013, outb => n1274);
   U1617 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_3_1_port, 
                           outb => n1013);
   U1618 : nand4 port map( a => n1280, b => n1281, c => n1282, d => n1283, outb
                           => n2290);
   U1619 : aoi22 port map( a => n1284, b => n1285, c => load_n_store_we_i, d =>
                           load_n_store_lazy_in_1_0_port, outb => n1283);
   U1620 : nor3 port map( a => n1286, b => n1287, c => n1288, outb => n1285);
   U1621 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_26_0_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_31_0_port, d =>
                           n370, outb => n1288);
   U1622 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_25_0_port, 
                           b => n507, outb => n1287);
   U1623 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_30_0_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_24_0_port, d =>
                           n509, outb => n1286);
   U1624 : nor3 port map( a => n1289, b => n1290, c => n512, outb => n1284);
   U1625 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_27_0_port, 
                           b => n513, outb => n1290);
   U1626 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_28_0_port,
                           b => n514, c => 
                           load_n_store_RGB_Array_1_block_ram_r_29_0_port, d =>
                           n515, outb => n1289);
   U1627 : nand4 port map( a => n516, b => n1291, c => n1292, d => n1293, outb 
                           => n1282);
   U1628 : nor3 port map( a => n1294, b => n1295, c => n1296, outb => n1293);
   U1629 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_18_0_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_23_0_port, d =>
                           n370, outb => n1296);
   U1630 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_17_0_port, 
                           b => n507, outb => n1295);
   U1631 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_22_0_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_16_0_port, d =>
                           n509, outb => n1294);
   U1632 : aoi22 port map( a => n523, b => n1297, c => n525, d => n1298, outb 
                           => n1292);
   U1633 : nand2 port map( a => n527, b => n1299, outb => n1291);
   U1634 : nand4 port map( a => n529, b => n1300, c => n1301, d => n1302, outb 
                           => n1281);
   U1635 : nor3 port map( a => n1303, b => n1304, c => n1305, outb => n1302);
   U1636 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_10_0_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_15_0_port, d =>
                           n370, outb => n1305);
   U1637 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_9_0_port, b
                           => n507, outb => n1304);
   U1638 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_14_0_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_8_0_port, d => 
                           n509, outb => n1303);
   U1639 : aoi22 port map( a => n523, b => n1306, c => n525, d => n1307, outb 
                           => n1301);
   U1640 : nand2 port map( a => n527, b => n950, outb => n1300);
   U1641 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_11_0_port,
                           outb => n950);
   U1642 : nand4 port map( a => n539, b => n1308, c => n1309, d => n1310, outb 
                           => n1280);
   U1643 : nor3 port map( a => n1311, b => n1312, c => n1313, outb => n1310);
   U1644 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_2_0_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_1_block_ram_r_7_0_port, d => 
                           n370, outb => n1313);
   U1645 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_1_0_port, b
                           => n507, outb => n1312);
   U1646 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_6_0_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_1_block_ram_r_0_0_port, d => 
                           n509, outb => n1311);
   U1647 : aoi22 port map( a => n523, b => n998, c => n525, d => n1006, outb =>
                           n1309);
   U1648 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_4_0_port, 
                           outb => n1006);
   U1649 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_5_0_port, 
                           outb => n998);
   U1650 : nand2 port map( a => n527, b => n1014, outb => n1308);
   U1651 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_3_0_port, 
                           outb => n1014);
   U1652 : oai22 port map( a => n199, b => n786, c => n787, d => n1314, outb =>
                           n2816);
   U1653 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_31_7_port,
                           outb => n1314);
   U1654 : oai22 port map( a => n197, b => n786, c => n787, d => n1315, outb =>
                           n2815);
   U1655 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_31_6_port,
                           outb => n1315);
   U1656 : oai22 port map( a => n195, b => n786, c => n787, d => n1316, outb =>
                           n2814);
   U1657 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_31_5_port,
                           outb => n1316);
   U1658 : oai22 port map( a => n193, b => n786, c => n787, d => n1317, outb =>
                           n2813);
   U1659 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_31_4_port,
                           outb => n1317);
   U1660 : oai22 port map( a => n191, b => n786, c => n787, d => n1318, outb =>
                           n2812);
   U1661 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_31_3_port,
                           outb => n1318);
   U1662 : oai22 port map( a => n189, b => n786, c => n787, d => n1319, outb =>
                           n2811);
   U1663 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_31_2_port,
                           outb => n1319);
   U1664 : oai22 port map( a => n187, b => n786, c => n787, d => n1320, outb =>
                           n2810);
   U1665 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_31_1_port,
                           outb => n1320);
   U1666 : oai22 port map( a => n185, b => n786, c => n787, d => n1321, outb =>
                           n2809);
   U1667 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_31_0_port,
                           outb => n1321);
   U1668 : oai22 port map( a => n199, b => n796, c => n797, d => n1322, outb =>
                           n2808);
   U1669 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_30_7_port,
                           outb => n1322);
   U1670 : oai22 port map( a => n197, b => n796, c => n797, d => n1323, outb =>
                           n2807);
   U1671 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_30_6_port,
                           outb => n1323);
   U1672 : oai22 port map( a => n195, b => n796, c => n797, d => n1324, outb =>
                           n2806);
   U1673 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_30_5_port,
                           outb => n1324);
   U1674 : oai22 port map( a => n193, b => n796, c => n797, d => n1325, outb =>
                           n2805);
   U1675 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_30_4_port,
                           outb => n1325);
   U1676 : oai22 port map( a => n191, b => n796, c => n797, d => n1326, outb =>
                           n2804);
   U1677 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_30_3_port,
                           outb => n1326);
   U1678 : oai22 port map( a => n189, b => n796, c => n797, d => n1327, outb =>
                           n2803);
   U1679 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_30_2_port,
                           outb => n1327);
   U1680 : oai22 port map( a => n187, b => n796, c => n797, d => n1328, outb =>
                           n2802);
   U1681 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_30_1_port,
                           outb => n1328);
   U1682 : oai22 port map( a => n185, b => n796, c => n797, d => n1329, outb =>
                           n2801);
   U1683 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_30_0_port,
                           outb => n1329);
   U1684 : oai22 port map( a => n199, b => n806, c => n807, d => n1330, outb =>
                           n2800);
   U1685 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_29_7_port,
                           outb => n1330);
   U1686 : oai22 port map( a => n197, b => n806, c => n807, d => n1331, outb =>
                           n2799);
   U1687 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_29_6_port,
                           outb => n1331);
   U1688 : oai22 port map( a => n195, b => n806, c => n807, d => n1332, outb =>
                           n2798);
   U1689 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_29_5_port,
                           outb => n1332);
   U1690 : oai22 port map( a => n193, b => n806, c => n807, d => n1333, outb =>
                           n2797);
   U1691 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_29_4_port,
                           outb => n1333);
   U1692 : oai22 port map( a => n191, b => n806, c => n807, d => n1334, outb =>
                           n2796);
   U1693 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_29_3_port,
                           outb => n1334);
   U1694 : oai22 port map( a => n189, b => n806, c => n807, d => n1335, outb =>
                           n2795);
   U1695 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_29_2_port,
                           outb => n1335);
   U1696 : oai22 port map( a => n187, b => n806, c => n807, d => n1336, outb =>
                           n2794);
   U1697 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_29_1_port,
                           outb => n1336);
   U1698 : oai22 port map( a => n185, b => n806, c => n807, d => n1337, outb =>
                           n2793);
   U1699 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_29_0_port,
                           outb => n1337);
   U1700 : oai22 port map( a => n199, b => n816, c => n817, d => n1338, outb =>
                           n2792);
   U1701 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_28_7_port,
                           outb => n1338);
   U1702 : oai22 port map( a => n197, b => n816, c => n817, d => n1339, outb =>
                           n2791);
   U1703 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_28_6_port,
                           outb => n1339);
   U1704 : oai22 port map( a => n195, b => n816, c => n817, d => n1340, outb =>
                           n2790);
   U1705 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_28_5_port,
                           outb => n1340);
   U1706 : oai22 port map( a => n193, b => n816, c => n817, d => n1341, outb =>
                           n2789);
   U1707 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_28_4_port,
                           outb => n1341);
   U1708 : oai22 port map( a => n191, b => n816, c => n817, d => n1342, outb =>
                           n2788);
   U1709 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_28_3_port,
                           outb => n1342);
   U1710 : oai22 port map( a => n189, b => n816, c => n817, d => n1343, outb =>
                           n2787);
   U1711 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_28_2_port,
                           outb => n1343);
   U1712 : oai22 port map( a => n187, b => n816, c => n817, d => n1344, outb =>
                           n2786);
   U1713 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_28_1_port,
                           outb => n1344);
   U1714 : oai22 port map( a => n185, b => n816, c => n817, d => n1345, outb =>
                           n2785);
   U1715 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_28_0_port,
                           outb => n1345);
   U1716 : oai22 port map( a => n199, b => n826, c => n827, d => n1346, outb =>
                           n2784);
   U1717 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_27_7_port,
                           outb => n1346);
   U1718 : oai22 port map( a => n197, b => n826, c => n827, d => n1347, outb =>
                           n2783);
   U1719 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_27_6_port,
                           outb => n1347);
   U1720 : oai22 port map( a => n195, b => n826, c => n827, d => n1348, outb =>
                           n2782);
   U1721 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_27_5_port,
                           outb => n1348);
   U1722 : oai22 port map( a => n193, b => n826, c => n827, d => n1349, outb =>
                           n2781);
   U1723 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_27_4_port,
                           outb => n1349);
   U1724 : oai22 port map( a => n191, b => n826, c => n827, d => n1350, outb =>
                           n2780);
   U1725 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_27_3_port,
                           outb => n1350);
   U1726 : oai22 port map( a => n189, b => n826, c => n827, d => n1351, outb =>
                           n2779);
   U1727 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_27_2_port,
                           outb => n1351);
   U1728 : oai22 port map( a => n187, b => n826, c => n827, d => n1352, outb =>
                           n2778);
   U1729 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_27_1_port,
                           outb => n1352);
   U1730 : oai22 port map( a => n185, b => n826, c => n827, d => n1353, outb =>
                           n2777);
   U1731 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_27_0_port,
                           outb => n1353);
   U1732 : oai22 port map( a => n199, b => n836, c => n837, d => n1354, outb =>
                           n2776);
   U1733 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_26_7_port,
                           outb => n1354);
   U1734 : oai22 port map( a => n197, b => n836, c => n837, d => n1355, outb =>
                           n2775);
   U1735 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_26_6_port,
                           outb => n1355);
   U1736 : oai22 port map( a => n195, b => n836, c => n837, d => n1356, outb =>
                           n2774);
   U1737 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_26_5_port,
                           outb => n1356);
   U1738 : oai22 port map( a => n193, b => n836, c => n837, d => n1357, outb =>
                           n2773);
   U1739 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_26_4_port,
                           outb => n1357);
   U1740 : oai22 port map( a => n191, b => n836, c => n837, d => n1358, outb =>
                           n2772);
   U1741 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_26_3_port,
                           outb => n1358);
   U1742 : oai22 port map( a => n189, b => n836, c => n837, d => n1359, outb =>
                           n2771);
   U1743 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_26_2_port,
                           outb => n1359);
   U1744 : oai22 port map( a => n187, b => n836, c => n837, d => n1360, outb =>
                           n2770);
   U1745 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_26_1_port,
                           outb => n1360);
   U1746 : oai22 port map( a => n185, b => n836, c => n837, d => n1361, outb =>
                           n2769);
   U1747 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_26_0_port,
                           outb => n1361);
   U1748 : oai22 port map( a => n199, b => n846, c => n847, d => n1362, outb =>
                           n2768);
   U1749 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_25_7_port,
                           outb => n1362);
   U1750 : oai22 port map( a => n197, b => n846, c => n847, d => n1363, outb =>
                           n2767);
   U1751 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_25_6_port,
                           outb => n1363);
   U1752 : oai22 port map( a => n195, b => n846, c => n847, d => n1364, outb =>
                           n2766);
   U1753 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_25_5_port,
                           outb => n1364);
   U1754 : oai22 port map( a => n193, b => n846, c => n847, d => n1365, outb =>
                           n2765);
   U1755 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_25_4_port,
                           outb => n1365);
   U1756 : oai22 port map( a => n191, b => n846, c => n847, d => n1366, outb =>
                           n2764);
   U1757 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_25_3_port,
                           outb => n1366);
   U1758 : oai22 port map( a => n189, b => n846, c => n847, d => n1367, outb =>
                           n2763);
   U1759 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_25_2_port,
                           outb => n1367);
   U1760 : oai22 port map( a => n187, b => n846, c => n847, d => n1368, outb =>
                           n2762);
   U1761 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_25_1_port,
                           outb => n1368);
   U1762 : oai22 port map( a => n185, b => n846, c => n847, d => n1369, outb =>
                           n2761);
   U1763 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_25_0_port,
                           outb => n1369);
   U1764 : oai22 port map( a => n199, b => n856, c => n857, d => n1370, outb =>
                           n2760);
   U1765 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_24_7_port,
                           outb => n1370);
   U1766 : oai22 port map( a => n197, b => n856, c => n857, d => n1371, outb =>
                           n2759);
   U1767 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_24_6_port,
                           outb => n1371);
   U1768 : oai22 port map( a => n195, b => n856, c => n857, d => n1372, outb =>
                           n2758);
   U1769 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_24_5_port,
                           outb => n1372);
   U1770 : oai22 port map( a => n193, b => n856, c => n857, d => n1373, outb =>
                           n2757);
   U1771 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_24_4_port,
                           outb => n1373);
   U1772 : oai22 port map( a => n191, b => n856, c => n857, d => n1374, outb =>
                           n2756);
   U1773 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_24_3_port,
                           outb => n1374);
   U1774 : oai22 port map( a => n189, b => n856, c => n857, d => n1375, outb =>
                           n2755);
   U1775 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_24_2_port,
                           outb => n1375);
   U1776 : oai22 port map( a => n187, b => n856, c => n857, d => n1376, outb =>
                           n2754);
   U1777 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_24_1_port,
                           outb => n1376);
   U1778 : oai22 port map( a => n185, b => n856, c => n857, d => n1377, outb =>
                           n2753);
   U1779 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_24_0_port,
                           outb => n1377);
   U1780 : oai22 port map( a => n199, b => n866, c => n867, d => n1378, outb =>
                           n2752);
   U1781 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_23_7_port,
                           outb => n1378);
   U1782 : oai22 port map( a => n197, b => n866, c => n867, d => n1379, outb =>
                           n2751);
   U1783 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_23_6_port,
                           outb => n1379);
   U1784 : oai22 port map( a => n195, b => n866, c => n867, d => n1380, outb =>
                           n2750);
   U1785 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_23_5_port,
                           outb => n1380);
   U1786 : oai22 port map( a => n193, b => n866, c => n867, d => n1381, outb =>
                           n2749);
   U1787 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_23_4_port,
                           outb => n1381);
   U1788 : oai22 port map( a => n191, b => n866, c => n867, d => n1382, outb =>
                           n2748);
   U1789 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_23_3_port,
                           outb => n1382);
   U1790 : oai22 port map( a => n189, b => n866, c => n867, d => n1383, outb =>
                           n2747);
   U1791 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_23_2_port,
                           outb => n1383);
   U1792 : oai22 port map( a => n187, b => n866, c => n867, d => n1384, outb =>
                           n2746);
   U1793 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_23_1_port,
                           outb => n1384);
   U1794 : oai22 port map( a => n185, b => n866, c => n867, d => n1385, outb =>
                           n2745);
   U1795 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_23_0_port,
                           outb => n1385);
   U1796 : oai22 port map( a => n199, b => n876, c => n877, d => n1386, outb =>
                           n2744);
   U1797 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_22_7_port,
                           outb => n1386);
   U1798 : oai22 port map( a => n197, b => n876, c => n877, d => n1387, outb =>
                           n2743);
   U1799 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_22_6_port,
                           outb => n1387);
   U1800 : oai22 port map( a => n195, b => n876, c => n877, d => n1388, outb =>
                           n2742);
   U1801 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_22_5_port,
                           outb => n1388);
   U1802 : oai22 port map( a => n193, b => n876, c => n877, d => n1389, outb =>
                           n2741);
   U1803 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_22_4_port,
                           outb => n1389);
   U1804 : oai22 port map( a => n191, b => n876, c => n877, d => n1390, outb =>
                           n2740);
   U1805 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_22_3_port,
                           outb => n1390);
   U1806 : oai22 port map( a => n189, b => n876, c => n877, d => n1391, outb =>
                           n2739);
   U1807 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_22_2_port,
                           outb => n1391);
   U1808 : oai22 port map( a => n187, b => n876, c => n877, d => n1392, outb =>
                           n2738);
   U1809 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_22_1_port,
                           outb => n1392);
   U1810 : oai22 port map( a => n185, b => n876, c => n877, d => n1393, outb =>
                           n2737);
   U1811 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_22_0_port,
                           outb => n1393);
   U1812 : oai22 port map( a => n199, b => n886, c => n887, d => n1056, outb =>
                           n2736);
   U1813 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_21_7_port,
                           outb => n1056);
   U1814 : oai22 port map( a => n197, b => n886, c => n887, d => n1091, outb =>
                           n2735);
   U1815 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_21_6_port,
                           outb => n1091);
   U1816 : oai22 port map( a => n195, b => n886, c => n887, d => n1126, outb =>
                           n2734);
   U1817 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_21_5_port,
                           outb => n1126);
   U1818 : oai22 port map( a => n193, b => n886, c => n887, d => n1161, outb =>
                           n2733);
   U1819 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_21_4_port,
                           outb => n1161);
   U1820 : oai22 port map( a => n191, b => n886, c => n887, d => n1195, outb =>
                           n2732);
   U1821 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_21_3_port,
                           outb => n1195);
   U1822 : oai22 port map( a => n189, b => n886, c => n887, d => n1229, outb =>
                           n2731);
   U1823 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_21_2_port,
                           outb => n1229);
   U1824 : oai22 port map( a => n187, b => n886, c => n887, d => n1263, outb =>
                           n2730);
   U1825 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_21_1_port,
                           outb => n1263);
   U1826 : oai22 port map( a => n185, b => n886, c => n887, d => n1297, outb =>
                           n2729);
   U1827 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_21_0_port,
                           outb => n1297);
   U1828 : oai22 port map( a => n199, b => n888, c => n889, d => n1057, outb =>
                           n2728);
   U1829 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_20_7_port,
                           outb => n1057);
   U1830 : oai22 port map( a => n197, b => n888, c => n889, d => n1092, outb =>
                           n2727);
   U1831 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_20_6_port,
                           outb => n1092);
   U1832 : oai22 port map( a => n195, b => n888, c => n889, d => n1127, outb =>
                           n2726);
   U1833 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_20_5_port,
                           outb => n1127);
   U1834 : oai22 port map( a => n193, b => n888, c => n889, d => n1162, outb =>
                           n2725);
   U1835 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_20_4_port,
                           outb => n1162);
   U1836 : oai22 port map( a => n191, b => n888, c => n889, d => n1196, outb =>
                           n2724);
   U1837 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_20_3_port,
                           outb => n1196);
   U1838 : oai22 port map( a => n189, b => n888, c => n889, d => n1230, outb =>
                           n2723);
   U1839 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_20_2_port,
                           outb => n1230);
   U1840 : oai22 port map( a => n187, b => n888, c => n889, d => n1264, outb =>
                           n2722);
   U1841 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_20_1_port,
                           outb => n1264);
   U1842 : oai22 port map( a => n185, b => n888, c => n889, d => n1298, outb =>
                           n2721);
   U1843 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_20_0_port,
                           outb => n1298);
   U1844 : oai22 port map( a => n199, b => n890, c => n891, d => n1058, outb =>
                           n2720);
   U1845 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_19_7_port,
                           outb => n1058);
   U1846 : oai22 port map( a => n197, b => n890, c => n891, d => n1093, outb =>
                           n2719);
   U1847 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_19_6_port,
                           outb => n1093);
   U1848 : oai22 port map( a => n195, b => n890, c => n891, d => n1128, outb =>
                           n2718);
   U1849 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_19_5_port,
                           outb => n1128);
   U1850 : oai22 port map( a => n193, b => n890, c => n891, d => n1163, outb =>
                           n2717);
   U1851 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_19_4_port,
                           outb => n1163);
   U1852 : oai22 port map( a => n191, b => n890, c => n891, d => n1197, outb =>
                           n2716);
   U1853 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_19_3_port,
                           outb => n1197);
   U1854 : oai22 port map( a => n189, b => n890, c => n891, d => n1231, outb =>
                           n2715);
   U1855 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_19_2_port,
                           outb => n1231);
   U1856 : oai22 port map( a => n187, b => n890, c => n891, d => n1265, outb =>
                           n2714);
   U1857 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_19_1_port,
                           outb => n1265);
   U1858 : oai22 port map( a => n185, b => n890, c => n891, d => n1299, outb =>
                           n2713);
   U1859 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_19_0_port,
                           outb => n1299);
   U1860 : oai22 port map( a => n199, b => n892, c => n893, d => n1394, outb =>
                           n2712);
   U1861 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_18_7_port,
                           outb => n1394);
   U1862 : oai22 port map( a => n197, b => n892, c => n893, d => n1395, outb =>
                           n2711);
   U1863 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_18_6_port,
                           outb => n1395);
   U1864 : oai22 port map( a => n195, b => n892, c => n893, d => n1396, outb =>
                           n2710);
   U1865 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_18_5_port,
                           outb => n1396);
   U1866 : oai22 port map( a => n193, b => n892, c => n893, d => n1397, outb =>
                           n2709);
   U1867 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_18_4_port,
                           outb => n1397);
   U1868 : oai22 port map( a => n191, b => n892, c => n893, d => n1398, outb =>
                           n2708);
   U1869 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_18_3_port,
                           outb => n1398);
   U1870 : oai22 port map( a => n189, b => n892, c => n893, d => n1399, outb =>
                           n2707);
   U1871 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_18_2_port,
                           outb => n1399);
   U1872 : oai22 port map( a => n187, b => n892, c => n893, d => n1400, outb =>
                           n2706);
   U1873 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_18_1_port,
                           outb => n1400);
   U1874 : oai22 port map( a => n185, b => n892, c => n893, d => n1401, outb =>
                           n2705);
   U1875 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_18_0_port,
                           outb => n1401);
   U1876 : oai22 port map( a => n199, b => n902, c => n903, d => n1402, outb =>
                           n2704);
   U1877 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_17_7_port,
                           outb => n1402);
   U1878 : oai22 port map( a => n197, b => n902, c => n903, d => n1403, outb =>
                           n2703);
   U1879 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_17_6_port,
                           outb => n1403);
   U1880 : oai22 port map( a => n195, b => n902, c => n903, d => n1404, outb =>
                           n2702);
   U1881 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_17_5_port,
                           outb => n1404);
   U1882 : oai22 port map( a => n193, b => n902, c => n903, d => n1405, outb =>
                           n2701);
   U1883 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_17_4_port,
                           outb => n1405);
   U1884 : oai22 port map( a => n191, b => n902, c => n903, d => n1406, outb =>
                           n2700);
   U1885 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_17_3_port,
                           outb => n1406);
   U1886 : oai22 port map( a => n189, b => n902, c => n903, d => n1407, outb =>
                           n2699);
   U1887 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_17_2_port,
                           outb => n1407);
   U1888 : oai22 port map( a => n187, b => n902, c => n903, d => n1408, outb =>
                           n2698);
   U1889 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_17_1_port,
                           outb => n1408);
   U1890 : oai22 port map( a => n185, b => n902, c => n903, d => n1409, outb =>
                           n2697);
   U1891 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_17_0_port,
                           outb => n1409);
   U1892 : oai22 port map( a => n199, b => n912, c => n913, d => n1410, outb =>
                           n2696);
   U1893 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_16_7_port,
                           outb => n1410);
   U1894 : oai22 port map( a => n197, b => n912, c => n913, d => n1411, outb =>
                           n2695);
   U1895 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_16_6_port,
                           outb => n1411);
   U1896 : oai22 port map( a => n195, b => n912, c => n913, d => n1412, outb =>
                           n2694);
   U1897 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_16_5_port,
                           outb => n1412);
   U1898 : oai22 port map( a => n193, b => n912, c => n913, d => n1413, outb =>
                           n2693);
   U1899 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_16_4_port,
                           outb => n1413);
   U1900 : oai22 port map( a => n191, b => n912, c => n913, d => n1414, outb =>
                           n2692);
   U1901 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_16_3_port,
                           outb => n1414);
   U1902 : oai22 port map( a => n189, b => n912, c => n913, d => n1415, outb =>
                           n2691);
   U1903 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_16_2_port,
                           outb => n1415);
   U1904 : oai22 port map( a => n187, b => n912, c => n913, d => n1416, outb =>
                           n2690);
   U1905 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_16_1_port,
                           outb => n1416);
   U1906 : oai22 port map( a => n185, b => n912, c => n913, d => n1417, outb =>
                           n2689);
   U1907 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_16_0_port,
                           outb => n1417);
   U1908 : oai22 port map( a => n199, b => n922, c => n923, d => n1418, outb =>
                           n2688);
   U1909 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_15_7_port,
                           outb => n1418);
   U1910 : oai22 port map( a => n197, b => n922, c => n923, d => n1419, outb =>
                           n2687);
   U1911 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_15_6_port,
                           outb => n1419);
   U1912 : oai22 port map( a => n195, b => n922, c => n923, d => n1420, outb =>
                           n2686);
   U1913 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_15_5_port,
                           outb => n1420);
   U1914 : oai22 port map( a => n193, b => n922, c => n923, d => n1421, outb =>
                           n2685);
   U1915 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_15_4_port,
                           outb => n1421);
   U1916 : oai22 port map( a => n191, b => n922, c => n923, d => n1422, outb =>
                           n2684);
   U1917 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_15_3_port,
                           outb => n1422);
   U1918 : oai22 port map( a => n189, b => n922, c => n923, d => n1423, outb =>
                           n2683);
   U1919 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_15_2_port,
                           outb => n1423);
   U1920 : oai22 port map( a => n187, b => n922, c => n923, d => n1424, outb =>
                           n2682);
   U1921 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_15_1_port,
                           outb => n1424);
   U1922 : oai22 port map( a => n185, b => n922, c => n923, d => n1425, outb =>
                           n2681);
   U1923 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_15_0_port,
                           outb => n1425);
   U1924 : oai22 port map( a => n199, b => n932, c => n933, d => n1426, outb =>
                           n2680);
   U1925 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_14_7_port,
                           outb => n1426);
   U1926 : oai22 port map( a => n197, b => n932, c => n933, d => n1427, outb =>
                           n2679);
   U1927 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_14_6_port,
                           outb => n1427);
   U1928 : oai22 port map( a => n195, b => n932, c => n933, d => n1428, outb =>
                           n2678);
   U1929 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_14_5_port,
                           outb => n1428);
   U1930 : oai22 port map( a => n193, b => n932, c => n933, d => n1429, outb =>
                           n2677);
   U1931 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_14_4_port,
                           outb => n1429);
   U1932 : oai22 port map( a => n191, b => n932, c => n933, d => n1430, outb =>
                           n2676);
   U1933 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_14_3_port,
                           outb => n1430);
   U1934 : oai22 port map( a => n189, b => n932, c => n933, d => n1431, outb =>
                           n2675);
   U1935 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_14_2_port,
                           outb => n1431);
   U1936 : oai22 port map( a => n187, b => n932, c => n933, d => n1432, outb =>
                           n2674);
   U1937 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_14_1_port,
                           outb => n1432);
   U1938 : oai22 port map( a => n185, b => n932, c => n933, d => n1433, outb =>
                           n2673);
   U1939 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_14_0_port,
                           outb => n1433);
   U1940 : oai22 port map( a => n199, b => n942, c => n943, d => n1065, outb =>
                           n2672);
   U1941 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_13_7_port,
                           outb => n1065);
   U1942 : oai22 port map( a => n197, b => n942, c => n943, d => n1100, outb =>
                           n2671);
   U1943 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_13_6_port,
                           outb => n1100);
   U1944 : oai22 port map( a => n195, b => n942, c => n943, d => n1135, outb =>
                           n2670);
   U1945 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_13_5_port,
                           outb => n1135);
   U1946 : oai22 port map( a => n193, b => n942, c => n943, d => n1170, outb =>
                           n2669);
   U1947 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_13_4_port,
                           outb => n1170);
   U1948 : oai22 port map( a => n191, b => n942, c => n943, d => n1204, outb =>
                           n2668);
   U1949 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_13_3_port,
                           outb => n1204);
   U1950 : oai22 port map( a => n189, b => n942, c => n943, d => n1238, outb =>
                           n2667);
   U1951 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_13_2_port,
                           outb => n1238);
   U1952 : oai22 port map( a => n187, b => n942, c => n943, d => n1272, outb =>
                           n2666);
   U1953 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_13_1_port,
                           outb => n1272);
   U1954 : oai22 port map( a => n185, b => n942, c => n943, d => n1306, outb =>
                           n2665);
   U1955 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_13_0_port,
                           outb => n1306);
   U1956 : oai22 port map( a => n199, b => n944, c => n945, d => n1066, outb =>
                           n2664);
   U1957 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_12_7_port,
                           outb => n1066);
   U1958 : oai22 port map( a => n197, b => n944, c => n945, d => n1101, outb =>
                           n2663);
   U1959 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_12_6_port,
                           outb => n1101);
   U1960 : oai22 port map( a => n195, b => n944, c => n945, d => n1136, outb =>
                           n2662);
   U1961 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_12_5_port,
                           outb => n1136);
   U1962 : oai22 port map( a => n193, b => n944, c => n945, d => n1171, outb =>
                           n2661);
   U1963 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_12_4_port,
                           outb => n1171);
   U1964 : inv port map( inb => load_n_store_lazy_in_1_4_port, outb => n193);
   U1965 : oai22 port map( a => n191, b => n944, c => n945, d => n1205, outb =>
                           n2660);
   U1966 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_12_3_port,
                           outb => n1205);
   U1967 : inv port map( inb => load_n_store_lazy_in_1_3_port, outb => n191);
   U1968 : oai22 port map( a => n189, b => n944, c => n945, d => n1239, outb =>
                           n2659);
   U1969 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_12_2_port,
                           outb => n1239);
   U1970 : inv port map( inb => load_n_store_lazy_in_1_2_port, outb => n189);
   U1971 : oai22 port map( a => n187, b => n944, c => n945, d => n1273, outb =>
                           n2658);
   U1972 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_12_1_port,
                           outb => n1273);
   U1973 : inv port map( inb => load_n_store_lazy_in_1_1_port, outb => n187);
   U1974 : oai22 port map( a => n185, b => n944, c => n945, d => n1307, outb =>
                           n2657);
   U1975 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_12_0_port,
                           outb => n1307);
   U1976 : inv port map( inb => load_n_store_lazy_in_1_0_port, outb => n185);
   U1977 : oai22 port map( a => n199, b => n380, c => n381, d => n1067, outb =>
                           n2656);
   U1978 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_11_7_port,
                           outb => n1067);
   U1979 : inv port map( inb => load_n_store_lazy_in_1_7_port, outb => n199);
   U1980 : oai22 port map( a => n197, b => n380, c => n381, d => n1102, outb =>
                           n2655);
   U1981 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_11_6_port,
                           outb => n1102);
   U1982 : inv port map( inb => load_n_store_lazy_in_1_6_port, outb => n197);
   U1983 : oai22 port map( a => n195, b => n380, c => n381, d => n1137, outb =>
                           n2654);
   U1984 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_11_5_port,
                           outb => n1137);
   U1985 : inv port map( inb => load_n_store_lazy_in_1_5_port, outb => n195);
   U1986 : oai22 port map( a => n209, b => n380, c => n381, d => n1434, outb =>
                           load_n_store_RGB_Array_0_n999);
   U1987 : oai22 port map( a => n207, b => n380, c => n381, d => n1435, outb =>
                           load_n_store_RGB_Array_0_n998);
   U1988 : oai22 port map( a => n205, b => n380, c => n381, d => n1436, outb =>
                           load_n_store_RGB_Array_0_n997);
   U1989 : oai22 port map( a => n203, b => n380, c => n381, d => n1437, outb =>
                           load_n_store_RGB_Array_0_n996);
   U1990 : oai22 port map( a => n201, b => n380, c => n381, d => n1438, outb =>
                           load_n_store_RGB_Array_0_n995);
   U1991 : oai22 port map( a => n215, b => n387, c => n388, d => n1439, outb =>
                           load_n_store_RGB_Array_0_n994);
   U1992 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_10_7_port,
                           outb => n1439);
   U1993 : oai22 port map( a => n213, b => n387, c => n388, d => n1440, outb =>
                           load_n_store_RGB_Array_0_n993);
   U1994 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_10_6_port,
                           outb => n1440);
   U1995 : oai22 port map( a => n211, b => n387, c => n388, d => n1441, outb =>
                           load_n_store_RGB_Array_0_n992);
   U1996 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_10_5_port,
                           outb => n1441);
   U1997 : oai22 port map( a => n209, b => n387, c => n388, d => n1442, outb =>
                           load_n_store_RGB_Array_0_n991);
   U1998 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_10_4_port,
                           outb => n1442);
   U1999 : oai22 port map( a => n207, b => n387, c => n388, d => n1443, outb =>
                           load_n_store_RGB_Array_0_n990);
   U2000 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_10_3_port,
                           outb => n1443);
   U2001 : oai22 port map( a => n205, b => n387, c => n388, d => n1444, outb =>
                           load_n_store_RGB_Array_0_n989);
   U2002 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_10_2_port,
                           outb => n1444);
   U2003 : oai22 port map( a => n203, b => n387, c => n388, d => n1445, outb =>
                           load_n_store_RGB_Array_0_n988);
   U2004 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_10_1_port,
                           outb => n1445);
   U2005 : oai22 port map( a => n201, b => n387, c => n388, d => n1446, outb =>
                           load_n_store_RGB_Array_0_n987);
   U2006 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_10_0_port,
                           outb => n1446);
   U2007 : inv port map( inb => n387, outb => n388);
   U2008 : nand2 port map( a => n1447, b => n1448, outb => n387);
   U2009 : oai22 port map( a => n215, b => n397, c => n398, d => n1449, outb =>
                           load_n_store_RGB_Array_0_n986);
   U2010 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_9_7_port, 
                           outb => n1449);
   U2011 : oai22 port map( a => n213, b => n397, c => n398, d => n1450, outb =>
                           load_n_store_RGB_Array_0_n985);
   U2012 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_9_6_port, 
                           outb => n1450);
   U2013 : oai22 port map( a => n211, b => n397, c => n398, d => n1451, outb =>
                           load_n_store_RGB_Array_0_n984);
   U2014 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_9_5_port, 
                           outb => n1451);
   U2015 : oai22 port map( a => n209, b => n397, c => n398, d => n1452, outb =>
                           load_n_store_RGB_Array_0_n983);
   U2016 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_9_4_port, 
                           outb => n1452);
   U2017 : oai22 port map( a => n207, b => n397, c => n398, d => n1453, outb =>
                           load_n_store_RGB_Array_0_n982);
   U2018 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_9_3_port, 
                           outb => n1453);
   U2019 : oai22 port map( a => n205, b => n397, c => n398, d => n1454, outb =>
                           load_n_store_RGB_Array_0_n981);
   U2020 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_9_2_port, 
                           outb => n1454);
   U2021 : oai22 port map( a => n203, b => n397, c => n398, d => n1455, outb =>
                           load_n_store_RGB_Array_0_n980);
   U2022 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_9_1_port, 
                           outb => n1455);
   U2023 : oai22 port map( a => n201, b => n397, c => n398, d => n1456, outb =>
                           load_n_store_RGB_Array_0_n979);
   U2024 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_9_0_port, 
                           outb => n1456);
   U2025 : inv port map( inb => n397, outb => n398);
   U2026 : nand2 port map( a => n1457, b => n1448, outb => n397);
   U2027 : oai22 port map( a => n215, b => n407, c => n408, d => n1458, outb =>
                           load_n_store_RGB_Array_0_n978);
   U2028 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_8_7_port, 
                           outb => n1458);
   U2029 : oai22 port map( a => n213, b => n407, c => n408, d => n1459, outb =>
                           load_n_store_RGB_Array_0_n977);
   U2030 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_8_6_port, 
                           outb => n1459);
   U2031 : oai22 port map( a => n211, b => n407, c => n408, d => n1460, outb =>
                           load_n_store_RGB_Array_0_n976);
   U2032 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_8_5_port, 
                           outb => n1460);
   U2033 : oai22 port map( a => n209, b => n407, c => n408, d => n1461, outb =>
                           load_n_store_RGB_Array_0_n975);
   U2034 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_8_4_port, 
                           outb => n1461);
   U2035 : oai22 port map( a => n207, b => n407, c => n408, d => n1462, outb =>
                           load_n_store_RGB_Array_0_n974);
   U2036 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_8_3_port, 
                           outb => n1462);
   U2037 : oai22 port map( a => n205, b => n407, c => n408, d => n1463, outb =>
                           load_n_store_RGB_Array_0_n973);
   U2038 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_8_2_port, 
                           outb => n1463);
   U2039 : oai22 port map( a => n203, b => n407, c => n408, d => n1464, outb =>
                           load_n_store_RGB_Array_0_n972);
   U2040 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_8_1_port, 
                           outb => n1464);
   U2041 : oai22 port map( a => n201, b => n407, c => n408, d => n1465, outb =>
                           load_n_store_RGB_Array_0_n971);
   U2042 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_8_0_port, 
                           outb => n1465);
   U2043 : inv port map( inb => n407, outb => n408);
   U2044 : nand2 port map( a => n1466, b => n1448, outb => n407);
   U2045 : oai22 port map( a => n215, b => n417, c => n418, d => n1467, outb =>
                           load_n_store_RGB_Array_0_n970);
   U2046 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_7_7_port, 
                           outb => n1467);
   U2047 : oai22 port map( a => n213, b => n417, c => n418, d => n1468, outb =>
                           load_n_store_RGB_Array_0_n969);
   U2048 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_7_6_port, 
                           outb => n1468);
   U2049 : oai22 port map( a => n211, b => n417, c => n418, d => n1469, outb =>
                           load_n_store_RGB_Array_0_n968);
   U2050 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_7_5_port, 
                           outb => n1469);
   U2051 : oai22 port map( a => n209, b => n417, c => n418, d => n1470, outb =>
                           load_n_store_RGB_Array_0_n967);
   U2052 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_7_4_port, 
                           outb => n1470);
   U2053 : oai22 port map( a => n207, b => n417, c => n418, d => n1471, outb =>
                           load_n_store_RGB_Array_0_n966);
   U2054 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_7_3_port, 
                           outb => n1471);
   U2055 : oai22 port map( a => n205, b => n417, c => n418, d => n1472, outb =>
                           load_n_store_RGB_Array_0_n965);
   U2056 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_7_2_port, 
                           outb => n1472);
   U2057 : oai22 port map( a => n203, b => n417, c => n418, d => n1473, outb =>
                           load_n_store_RGB_Array_0_n964);
   U2058 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_7_1_port, 
                           outb => n1473);
   U2059 : oai22 port map( a => n201, b => n417, c => n418, d => n1474, outb =>
                           load_n_store_RGB_Array_0_n963);
   U2060 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_7_0_port, 
                           outb => n1474);
   U2061 : inv port map( inb => n417, outb => n418);
   U2062 : nand2 port map( a => n1475, b => n1476, outb => n417);
   U2063 : oai22 port map( a => n215, b => n427, c => n428, d => n1477, outb =>
                           load_n_store_RGB_Array_0_n962);
   U2064 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_6_7_port, 
                           outb => n1477);
   U2065 : oai22 port map( a => n213, b => n427, c => n428, d => n1478, outb =>
                           load_n_store_RGB_Array_0_n961);
   U2066 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_6_6_port, 
                           outb => n1478);
   U2067 : oai22 port map( a => n211, b => n427, c => n428, d => n1479, outb =>
                           load_n_store_RGB_Array_0_n960);
   U2068 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_6_5_port, 
                           outb => n1479);
   U2069 : oai22 port map( a => n209, b => n427, c => n428, d => n1480, outb =>
                           load_n_store_RGB_Array_0_n959);
   U2070 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_6_4_port, 
                           outb => n1480);
   U2071 : oai22 port map( a => n207, b => n427, c => n428, d => n1481, outb =>
                           load_n_store_RGB_Array_0_n958);
   U2072 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_6_3_port, 
                           outb => n1481);
   U2073 : oai22 port map( a => n205, b => n427, c => n428, d => n1482, outb =>
                           load_n_store_RGB_Array_0_n957);
   U2074 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_6_2_port, 
                           outb => n1482);
   U2075 : oai22 port map( a => n203, b => n427, c => n428, d => n1483, outb =>
                           load_n_store_RGB_Array_0_n956);
   U2076 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_6_1_port, 
                           outb => n1483);
   U2077 : oai22 port map( a => n201, b => n427, c => n428, d => n1484, outb =>
                           load_n_store_RGB_Array_0_n955);
   U2078 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_6_0_port, 
                           outb => n1484);
   U2079 : inv port map( inb => n427, outb => n428);
   U2080 : nand2 port map( a => n1485, b => n1475, outb => n427);
   U2081 : oai22 port map( a => n215, b => n437, c => n438, d => n1486, outb =>
                           load_n_store_RGB_Array_0_n954);
   U2082 : oai22 port map( a => n213, b => n437, c => n438, d => n1487, outb =>
                           load_n_store_RGB_Array_0_n953);
   U2083 : oai22 port map( a => n211, b => n437, c => n438, d => n1488, outb =>
                           load_n_store_RGB_Array_0_n952);
   U2084 : oai22 port map( a => n209, b => n437, c => n438, d => n1489, outb =>
                           load_n_store_RGB_Array_0_n951);
   U2085 : oai22 port map( a => n207, b => n437, c => n438, d => n1490, outb =>
                           load_n_store_RGB_Array_0_n950);
   U2086 : oai22 port map( a => n205, b => n437, c => n438, d => n1491, outb =>
                           load_n_store_RGB_Array_0_n949);
   U2087 : oai22 port map( a => n203, b => n437, c => n438, d => n1492, outb =>
                           load_n_store_RGB_Array_0_n948);
   U2088 : oai22 port map( a => n201, b => n437, c => n438, d => n1493, outb =>
                           load_n_store_RGB_Array_0_n947);
   U2089 : inv port map( inb => n437, outb => n438);
   U2090 : nand2 port map( a => n523, b => n1475, outb => n437);
   U2091 : oai22 port map( a => n215, b => n447, c => n448, d => n1494, outb =>
                           load_n_store_RGB_Array_0_n946);
   U2092 : oai22 port map( a => n213, b => n447, c => n448, d => n1495, outb =>
                           load_n_store_RGB_Array_0_n945);
   U2093 : oai22 port map( a => n211, b => n447, c => n448, d => n1496, outb =>
                           load_n_store_RGB_Array_0_n944);
   U2094 : oai22 port map( a => n209, b => n447, c => n448, d => n1497, outb =>
                           load_n_store_RGB_Array_0_n943);
   U2095 : oai22 port map( a => n207, b => n447, c => n448, d => n1498, outb =>
                           load_n_store_RGB_Array_0_n942);
   U2096 : oai22 port map( a => n205, b => n447, c => n448, d => n1499, outb =>
                           load_n_store_RGB_Array_0_n941);
   U2097 : oai22 port map( a => n203, b => n447, c => n448, d => n1500, outb =>
                           load_n_store_RGB_Array_0_n940);
   U2098 : oai22 port map( a => n201, b => n447, c => n448, d => n1501, outb =>
                           load_n_store_RGB_Array_0_n939);
   U2099 : inv port map( inb => n447, outb => n448);
   U2100 : nand2 port map( a => n525, b => n1475, outb => n447);
   U2101 : oai22 port map( a => n215, b => n457, c => n458, d => n1502, outb =>
                           load_n_store_RGB_Array_0_n938);
   U2102 : oai22 port map( a => n213, b => n457, c => n458, d => n1503, outb =>
                           load_n_store_RGB_Array_0_n937);
   U2103 : oai22 port map( a => n211, b => n457, c => n458, d => n1504, outb =>
                           load_n_store_RGB_Array_0_n936);
   U2104 : oai22 port map( a => n209, b => n457, c => n458, d => n1505, outb =>
                           load_n_store_RGB_Array_0_n935);
   U2105 : oai22 port map( a => n207, b => n457, c => n458, d => n1506, outb =>
                           load_n_store_RGB_Array_0_n934);
   U2106 : oai22 port map( a => n205, b => n457, c => n458, d => n1507, outb =>
                           load_n_store_RGB_Array_0_n933);
   U2107 : oai22 port map( a => n203, b => n457, c => n458, d => n1508, outb =>
                           load_n_store_RGB_Array_0_n932);
   U2108 : oai22 port map( a => n201, b => n457, c => n458, d => n1509, outb =>
                           load_n_store_RGB_Array_0_n931);
   U2109 : inv port map( inb => n457, outb => n458);
   U2110 : nand2 port map( a => n1475, b => n527, outb => n457);
   U2111 : oai22 port map( a => n215, b => n467, c => n468, d => n1510, outb =>
                           load_n_store_RGB_Array_0_n930);
   U2112 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_2_7_port, 
                           outb => n1510);
   U2113 : oai22 port map( a => n213, b => n467, c => n468, d => n1511, outb =>
                           load_n_store_RGB_Array_0_n929);
   U2114 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_2_6_port, 
                           outb => n1511);
   U2115 : oai22 port map( a => n211, b => n467, c => n468, d => n1512, outb =>
                           load_n_store_RGB_Array_0_n928);
   U2116 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_2_5_port, 
                           outb => n1512);
   U2117 : oai22 port map( a => n209, b => n467, c => n468, d => n1513, outb =>
                           load_n_store_RGB_Array_0_n927);
   U2118 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_2_4_port, 
                           outb => n1513);
   U2119 : oai22 port map( a => n207, b => n467, c => n468, d => n1514, outb =>
                           load_n_store_RGB_Array_0_n926);
   U2120 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_2_3_port, 
                           outb => n1514);
   U2121 : oai22 port map( a => n205, b => n467, c => n468, d => n1515, outb =>
                           load_n_store_RGB_Array_0_n925);
   U2122 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_2_2_port, 
                           outb => n1515);
   U2123 : oai22 port map( a => n203, b => n467, c => n468, d => n1516, outb =>
                           load_n_store_RGB_Array_0_n924);
   U2124 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_2_1_port, 
                           outb => n1516);
   U2125 : oai22 port map( a => n201, b => n467, c => n468, d => n1517, outb =>
                           load_n_store_RGB_Array_0_n923);
   U2126 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_2_0_port, 
                           outb => n1517);
   U2127 : inv port map( inb => n467, outb => n468);
   U2128 : nand2 port map( a => n1475, b => n1447, outb => n467);
   U2129 : oai22 port map( a => n215, b => n477, c => n478, d => n1518, outb =>
                           load_n_store_RGB_Array_0_n922);
   U2130 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_1_7_port, 
                           outb => n1518);
   U2131 : oai22 port map( a => n213, b => n477, c => n478, d => n1519, outb =>
                           load_n_store_RGB_Array_0_n921);
   U2132 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_1_6_port, 
                           outb => n1519);
   U2133 : oai22 port map( a => n211, b => n477, c => n478, d => n1520, outb =>
                           load_n_store_RGB_Array_0_n920);
   U2134 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_1_5_port, 
                           outb => n1520);
   U2135 : oai22 port map( a => n209, b => n477, c => n478, d => n1521, outb =>
                           load_n_store_RGB_Array_0_n919);
   U2136 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_1_4_port, 
                           outb => n1521);
   U2137 : oai22 port map( a => n207, b => n477, c => n478, d => n1522, outb =>
                           load_n_store_RGB_Array_0_n918);
   U2138 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_1_3_port, 
                           outb => n1522);
   U2139 : oai22 port map( a => n205, b => n477, c => n478, d => n1523, outb =>
                           load_n_store_RGB_Array_0_n917);
   U2140 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_1_2_port, 
                           outb => n1523);
   U2141 : oai22 port map( a => n203, b => n477, c => n478, d => n1524, outb =>
                           load_n_store_RGB_Array_0_n916);
   U2142 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_1_1_port, 
                           outb => n1524);
   U2143 : oai22 port map( a => n201, b => n477, c => n478, d => n1525, outb =>
                           load_n_store_RGB_Array_0_n915);
   U2144 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_1_0_port, 
                           outb => n1525);
   U2145 : inv port map( inb => n477, outb => n478);
   U2146 : nand2 port map( a => n1475, b => n1457, outb => n477);
   U2147 : oai22 port map( a => n215, b => n487, c => n488, d => n1526, outb =>
                           load_n_store_RGB_Array_0_n914);
   U2148 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_0_7_port, 
                           outb => n1526);
   U2149 : oai22 port map( a => n213, b => n487, c => n488, d => n1527, outb =>
                           load_n_store_RGB_Array_0_n913);
   U2150 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_0_6_port, 
                           outb => n1527);
   U2151 : oai22 port map( a => n211, b => n487, c => n488, d => n1528, outb =>
                           load_n_store_RGB_Array_0_n912);
   U2152 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_0_5_port, 
                           outb => n1528);
   U2153 : oai22 port map( a => n209, b => n487, c => n488, d => n1529, outb =>
                           load_n_store_RGB_Array_0_n911);
   U2154 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_0_4_port, 
                           outb => n1529);
   U2155 : oai22 port map( a => n207, b => n487, c => n488, d => n1530, outb =>
                           load_n_store_RGB_Array_0_n910);
   U2156 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_0_3_port, 
                           outb => n1530);
   U2157 : oai22 port map( a => n205, b => n487, c => n488, d => n1531, outb =>
                           load_n_store_RGB_Array_0_n909);
   U2158 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_0_2_port, 
                           outb => n1531);
   U2159 : oai22 port map( a => n203, b => n487, c => n488, d => n1532, outb =>
                           load_n_store_RGB_Array_0_n908);
   U2160 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_0_1_port, 
                           outb => n1532);
   U2161 : oai22 port map( a => n201, b => n487, c => n488, d => n1533, outb =>
                           load_n_store_RGB_Array_0_n907);
   U2162 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_0_0_port, 
                           outb => n1533);
   U2163 : inv port map( inb => n487, outb => n488);
   U2164 : nand2 port map( a => n1475, b => n1466, outb => n487);
   U2165 : nor3 port map( a => load_n_store_s_addr_3_port, b => 
                           load_n_store_s_addr_4_port, c => n1534, outb => 
                           n1475);
   U2166 : nand4 port map( a => n1535, b => n1536, c => n1537, d => n1538, outb
                           => load_n_store_RGB_Array_0_n657);
   U2167 : aoi22 port map( a => n1539, b => n1540, c => load_n_store_we_i, d =>
                           load_n_store_lazy_in_0_7_port, outb => n1538);
   U2168 : nor3 port map( a => n1541, b => n1542, c => n1543, outb => n1540);
   U2169 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_26_7_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_31_7_port, d =>
                           n370, outb => n1543);
   U2170 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_25_7_port, 
                           b => n507, outb => n1542);
   U2171 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_30_7_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_24_7_port, d =>
                           n509, outb => n1541);
   U2172 : nor3 port map( a => n1544, b => n1545, c => n512, outb => n1539);
   U2173 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_27_7_port, 
                           b => n513, outb => n1545);
   U2174 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_28_7_port,
                           b => n514, c => 
                           load_n_store_RGB_Array_0_block_ram_r_29_7_port, d =>
                           n515, outb => n1544);
   U2175 : nand4 port map( a => n516, b => n1546, c => n1547, d => n1548, outb 
                           => n1537);
   U2176 : nor3 port map( a => n1549, b => n1550, c => n1551, outb => n1548);
   U2177 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_18_7_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_23_7_port, d =>
                           n370, outb => n1551);
   U2178 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_17_7_port, 
                           b => n507, outb => n1550);
   U2179 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_22_7_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_16_7_port, d =>
                           n509, outb => n1549);
   U2180 : aoi22 port map( a => n523, b => n1552, c => n525, d => n1553, outb 
                           => n1547);
   U2181 : nand2 port map( a => n527, b => n1554, outb => n1546);
   U2182 : nand4 port map( a => n529, b => n1555, c => n1556, d => n1557, outb 
                           => n1536);
   U2183 : nor3 port map( a => n1558, b => n1559, c => n1560, outb => n1557);
   U2184 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_10_7_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_15_7_port, d =>
                           n370, outb => n1560);
   U2185 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_9_7_port, b
                           => n507, outb => n1559);
   U2186 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_14_7_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_8_7_port, d => 
                           n509, outb => n1558);
   U2187 : aoi22 port map( a => n523, b => n1561, c => n525, d => n1562, outb 
                           => n1556);
   U2188 : nand2 port map( a => n527, b => n1563, outb => n1555);
   U2189 : nand4 port map( a => n539, b => n1564, c => n1565, d => n1566, outb 
                           => n1535);
   U2190 : nor3 port map( a => n1567, b => n1568, c => n1569, outb => n1566);
   U2191 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_2_7_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_7_7_port, d => 
                           n370, outb => n1569);
   U2192 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_1_7_port, b
                           => n507, outb => n1568);
   U2193 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_6_7_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_0_7_port, d => 
                           n509, outb => n1567);
   U2194 : aoi22 port map( a => n523, b => n1486, c => n525, d => n1494, outb 
                           => n1565);
   U2195 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_4_7_port, 
                           outb => n1494);
   U2196 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_5_7_port, 
                           outb => n1486);
   U2197 : nand2 port map( a => n527, b => n1502, outb => n1564);
   U2198 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_3_7_port, 
                           outb => n1502);
   U2199 : nand4 port map( a => n1570, b => n1571, c => n1572, d => n1573, outb
                           => load_n_store_RGB_Array_0_n654);
   U2200 : aoi22 port map( a => n1574, b => n1575, c => load_n_store_we_i, d =>
                           load_n_store_lazy_in_0_6_port, outb => n1573);
   U2201 : nor3 port map( a => n1576, b => n1577, c => n1578, outb => n1575);
   U2202 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_26_6_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_31_6_port, d =>
                           n370, outb => n1578);
   U2203 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_25_6_port, 
                           b => n507, outb => n1577);
   U2204 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_30_6_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_24_6_port, d =>
                           n509, outb => n1576);
   U2205 : nor3 port map( a => n1579, b => n1580, c => n512, outb => n1574);
   U2206 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_27_6_port, 
                           b => n513, outb => n1580);
   U2207 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_28_6_port,
                           b => n514, c => 
                           load_n_store_RGB_Array_0_block_ram_r_29_6_port, d =>
                           n515, outb => n1579);
   U2208 : nand4 port map( a => n516, b => n1581, c => n1582, d => n1583, outb 
                           => n1572);
   U2209 : nor3 port map( a => n1584, b => n1585, c => n1586, outb => n1583);
   U2210 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_18_6_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_23_6_port, d =>
                           n370, outb => n1586);
   U2211 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_17_6_port, 
                           b => n507, outb => n1585);
   U2212 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_22_6_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_16_6_port, d =>
                           n509, outb => n1584);
   U2213 : aoi22 port map( a => n523, b => n1587, c => n525, d => n1588, outb 
                           => n1582);
   U2214 : nand2 port map( a => n527, b => n1589, outb => n1581);
   U2215 : nand4 port map( a => n529, b => n1590, c => n1591, d => n1592, outb 
                           => n1571);
   U2216 : nor3 port map( a => n1593, b => n1594, c => n1595, outb => n1592);
   U2217 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_10_6_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_15_6_port, d =>
                           n370, outb => n1595);
   U2218 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_9_6_port, b
                           => n507, outb => n1594);
   U2219 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_14_6_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_8_6_port, d => 
                           n509, outb => n1593);
   U2220 : aoi22 port map( a => n523, b => n1596, c => n525, d => n1597, outb 
                           => n1591);
   U2221 : nand2 port map( a => n527, b => n1598, outb => n1590);
   U2222 : nand4 port map( a => n539, b => n1599, c => n1600, d => n1601, outb 
                           => n1570);
   U2223 : nor3 port map( a => n1602, b => n1603, c => n1604, outb => n1601);
   U2224 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_2_6_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_7_6_port, d => 
                           n370, outb => n1604);
   U2225 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_1_6_port, b
                           => n507, outb => n1603);
   U2226 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_6_6_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_0_6_port, d => 
                           n509, outb => n1602);
   U2227 : aoi22 port map( a => n523, b => n1487, c => n525, d => n1495, outb 
                           => n1600);
   U2228 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_4_6_port, 
                           outb => n1495);
   U2229 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_5_6_port, 
                           outb => n1487);
   U2230 : nand2 port map( a => n527, b => n1503, outb => n1599);
   U2231 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_3_6_port, 
                           outb => n1503);
   U2232 : nand4 port map( a => n1605, b => n1606, c => n1607, d => n1608, outb
                           => load_n_store_RGB_Array_0_n651);
   U2233 : aoi22 port map( a => n1609, b => n1610, c => load_n_store_we_i, d =>
                           load_n_store_lazy_in_0_5_port, outb => n1608);
   U2234 : nor3 port map( a => n1611, b => n1612, c => n1613, outb => n1610);
   U2235 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_26_5_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_31_5_port, d =>
                           n370, outb => n1613);
   U2236 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_25_5_port, 
                           b => n507, outb => n1612);
   U2237 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_30_5_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_24_5_port, d =>
                           n509, outb => n1611);
   U2238 : nor3 port map( a => n1614, b => n1615, c => n512, outb => n1609);
   U2239 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_27_5_port, 
                           b => n513, outb => n1615);
   U2240 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_28_5_port,
                           b => n514, c => 
                           load_n_store_RGB_Array_0_block_ram_r_29_5_port, d =>
                           n515, outb => n1614);
   U2241 : nand4 port map( a => n516, b => n1616, c => n1617, d => n1618, outb 
                           => n1607);
   U2242 : nor3 port map( a => n1619, b => n1620, c => n1621, outb => n1618);
   U2243 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_18_5_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_23_5_port, d =>
                           n370, outb => n1621);
   U2244 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_17_5_port, 
                           b => n507, outb => n1620);
   U2245 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_22_5_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_16_5_port, d =>
                           n509, outb => n1619);
   U2246 : aoi22 port map( a => n523, b => n1622, c => n525, d => n1623, outb 
                           => n1617);
   U2247 : nand2 port map( a => n527, b => n1624, outb => n1616);
   U2248 : nand4 port map( a => n529, b => n1625, c => n1626, d => n1627, outb 
                           => n1606);
   U2249 : nor3 port map( a => n1628, b => n1629, c => n1630, outb => n1627);
   U2250 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_10_5_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_15_5_port, d =>
                           n370, outb => n1630);
   U2251 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_9_5_port, b
                           => n507, outb => n1629);
   U2252 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_14_5_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_8_5_port, d => 
                           n509, outb => n1628);
   U2253 : aoi22 port map( a => n523, b => n1631, c => n525, d => n1632, outb 
                           => n1626);
   U2254 : nand2 port map( a => n527, b => n1633, outb => n1625);
   U2255 : nand4 port map( a => n539, b => n1634, c => n1635, d => n1636, outb 
                           => n1605);
   U2256 : nor3 port map( a => n1637, b => n1638, c => n1639, outb => n1636);
   U2257 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_2_5_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_7_5_port, d => 
                           n370, outb => n1639);
   U2258 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_1_5_port, b
                           => n507, outb => n1638);
   U2259 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_6_5_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_0_5_port, d => 
                           n509, outb => n1637);
   U2260 : aoi22 port map( a => n523, b => n1488, c => n525, d => n1496, outb 
                           => n1635);
   U2261 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_4_5_port, 
                           outb => n1496);
   U2262 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_5_5_port, 
                           outb => n1488);
   U2263 : nand2 port map( a => n527, b => n1504, outb => n1634);
   U2264 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_3_5_port, 
                           outb => n1504);
   U2265 : nand4 port map( a => n1640, b => n1641, c => n1642, d => n1643, outb
                           => load_n_store_RGB_Array_0_n648);
   U2266 : aoi22 port map( a => n1644, b => n1645, c => load_n_store_we_i, d =>
                           load_n_store_lazy_in_0_4_port, outb => n1643);
   U2267 : nor3 port map( a => n1646, b => n1647, c => n1648, outb => n1645);
   U2268 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_26_4_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_31_4_port, d =>
                           n370, outb => n1648);
   U2269 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_25_4_port, 
                           b => n507, outb => n1647);
   U2270 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_30_4_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_24_4_port, d =>
                           n509, outb => n1646);
   U2271 : nor3 port map( a => n1649, b => n1650, c => n512, outb => n1644);
   U2272 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_27_4_port, 
                           b => n513, outb => n1650);
   U2273 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_28_4_port,
                           b => n514, c => 
                           load_n_store_RGB_Array_0_block_ram_r_29_4_port, d =>
                           n515, outb => n1649);
   U2274 : nand4 port map( a => n516, b => n1651, c => n1652, d => n1653, outb 
                           => n1642);
   U2275 : nor3 port map( a => n1654, b => n1655, c => n1656, outb => n1653);
   U2276 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_18_4_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_23_4_port, d =>
                           n370, outb => n1656);
   U2277 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_17_4_port, 
                           b => n507, outb => n1655);
   U2278 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_22_4_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_16_4_port, d =>
                           n509, outb => n1654);
   U2279 : aoi22 port map( a => n523, b => n1657, c => n525, d => n1658, outb 
                           => n1652);
   U2280 : nand2 port map( a => n527, b => n1659, outb => n1651);
   U2281 : nand4 port map( a => n529, b => n1660, c => n1661, d => n1662, outb 
                           => n1641);
   U2282 : nor3 port map( a => n1663, b => n1664, c => n1665, outb => n1662);
   U2283 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_10_4_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_15_4_port, d =>
                           n370, outb => n1665);
   U2284 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_9_4_port, b
                           => n507, outb => n1664);
   U2285 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_14_4_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_8_4_port, d => 
                           n509, outb => n1663);
   U2286 : aoi22 port map( a => n523, b => n1666, c => n525, d => n1667, outb 
                           => n1661);
   U2287 : nand2 port map( a => n527, b => n1434, outb => n1660);
   U2288 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_11_4_port,
                           outb => n1434);
   U2289 : nand4 port map( a => n539, b => n1668, c => n1669, d => n1670, outb 
                           => n1640);
   U2290 : nor3 port map( a => n1671, b => n1672, c => n1673, outb => n1670);
   U2291 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_2_4_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_7_4_port, d => 
                           n370, outb => n1673);
   U2292 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_1_4_port, b
                           => n507, outb => n1672);
   U2293 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_6_4_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_0_4_port, d => 
                           n509, outb => n1671);
   U2294 : aoi22 port map( a => n523, b => n1489, c => n525, d => n1497, outb 
                           => n1669);
   U2295 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_4_4_port, 
                           outb => n1497);
   U2296 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_5_4_port, 
                           outb => n1489);
   U2297 : nand2 port map( a => n527, b => n1505, outb => n1668);
   U2298 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_3_4_port, 
                           outb => n1505);
   U2299 : nand4 port map( a => n1674, b => n1675, c => n1676, d => n1677, outb
                           => load_n_store_RGB_Array_0_n645);
   U2300 : aoi22 port map( a => n1678, b => n1679, c => load_n_store_we_i, d =>
                           load_n_store_lazy_in_0_3_port, outb => n1677);
   U2301 : nor3 port map( a => n1680, b => n1681, c => n1682, outb => n1679);
   U2302 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_26_3_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_31_3_port, d =>
                           n370, outb => n1682);
   U2303 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_25_3_port, 
                           b => n507, outb => n1681);
   U2304 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_30_3_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_24_3_port, d =>
                           n509, outb => n1680);
   U2305 : nor3 port map( a => n1683, b => n1684, c => n512, outb => n1678);
   U2306 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_27_3_port, 
                           b => n513, outb => n1684);
   U2307 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_28_3_port,
                           b => n514, c => 
                           load_n_store_RGB_Array_0_block_ram_r_29_3_port, d =>
                           n515, outb => n1683);
   U2308 : nand4 port map( a => n516, b => n1685, c => n1686, d => n1687, outb 
                           => n1676);
   U2309 : nor3 port map( a => n1688, b => n1689, c => n1690, outb => n1687);
   U2310 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_18_3_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_23_3_port, d =>
                           n370, outb => n1690);
   U2311 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_17_3_port, 
                           b => n507, outb => n1689);
   U2312 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_22_3_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_16_3_port, d =>
                           n509, outb => n1688);
   U2313 : aoi22 port map( a => n523, b => n1691, c => n525, d => n1692, outb 
                           => n1686);
   U2314 : nand2 port map( a => n527, b => n1693, outb => n1685);
   U2315 : nand4 port map( a => n529, b => n1694, c => n1695, d => n1696, outb 
                           => n1675);
   U2316 : nor3 port map( a => n1697, b => n1698, c => n1699, outb => n1696);
   U2317 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_10_3_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_15_3_port, d =>
                           n370, outb => n1699);
   U2318 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_9_3_port, b
                           => n507, outb => n1698);
   U2319 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_14_3_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_8_3_port, d => 
                           n509, outb => n1697);
   U2320 : aoi22 port map( a => n523, b => n1700, c => n525, d => n1701, outb 
                           => n1695);
   U2321 : nand2 port map( a => n527, b => n1435, outb => n1694);
   U2322 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_11_3_port,
                           outb => n1435);
   U2323 : nand4 port map( a => n539, b => n1702, c => n1703, d => n1704, outb 
                           => n1674);
   U2324 : nor3 port map( a => n1705, b => n1706, c => n1707, outb => n1704);
   U2325 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_2_3_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_7_3_port, d => 
                           n370, outb => n1707);
   U2326 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_1_3_port, b
                           => n507, outb => n1706);
   U2327 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_6_3_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_0_3_port, d => 
                           n509, outb => n1705);
   U2328 : aoi22 port map( a => n523, b => n1490, c => n525, d => n1498, outb 
                           => n1703);
   U2329 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_4_3_port, 
                           outb => n1498);
   U2330 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_5_3_port, 
                           outb => n1490);
   U2331 : nand2 port map( a => n527, b => n1506, outb => n1702);
   U2332 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_3_3_port, 
                           outb => n1506);
   U2333 : nand4 port map( a => n1708, b => n1709, c => n1710, d => n1711, outb
                           => load_n_store_RGB_Array_0_n642);
   U2334 : aoi22 port map( a => n1712, b => n1713, c => load_n_store_we_i, d =>
                           load_n_store_lazy_in_0_2_port, outb => n1711);
   U2335 : nor3 port map( a => n1714, b => n1715, c => n1716, outb => n1713);
   U2336 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_26_2_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_31_2_port, d =>
                           n370, outb => n1716);
   U2337 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_25_2_port, 
                           b => n507, outb => n1715);
   U2338 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_30_2_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_24_2_port, d =>
                           n509, outb => n1714);
   U2339 : nor3 port map( a => n1717, b => n1718, c => n512, outb => n1712);
   U2340 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_27_2_port, 
                           b => n513, outb => n1718);
   U2341 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_28_2_port,
                           b => n514, c => 
                           load_n_store_RGB_Array_0_block_ram_r_29_2_port, d =>
                           n515, outb => n1717);
   U2342 : nand4 port map( a => n516, b => n1719, c => n1720, d => n1721, outb 
                           => n1710);
   U2343 : nor3 port map( a => n1722, b => n1723, c => n1724, outb => n1721);
   U2344 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_18_2_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_23_2_port, d =>
                           n370, outb => n1724);
   U2345 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_17_2_port, 
                           b => n507, outb => n1723);
   U2346 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_22_2_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_16_2_port, d =>
                           n509, outb => n1722);
   U2347 : aoi22 port map( a => n523, b => n1725, c => n525, d => n1726, outb 
                           => n1720);
   U2348 : nand2 port map( a => n527, b => n1727, outb => n1719);
   U2349 : nand4 port map( a => n529, b => n1728, c => n1729, d => n1730, outb 
                           => n1709);
   U2350 : nor3 port map( a => n1731, b => n1732, c => n1733, outb => n1730);
   U2351 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_10_2_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_15_2_port, d =>
                           n370, outb => n1733);
   U2352 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_9_2_port, b
                           => n507, outb => n1732);
   U2353 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_14_2_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_8_2_port, d => 
                           n509, outb => n1731);
   U2354 : aoi22 port map( a => n523, b => n1734, c => n525, d => n1735, outb 
                           => n1729);
   U2355 : nand2 port map( a => n527, b => n1436, outb => n1728);
   U2356 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_11_2_port,
                           outb => n1436);
   U2357 : nand4 port map( a => n539, b => n1736, c => n1737, d => n1738, outb 
                           => n1708);
   U2358 : nor3 port map( a => n1739, b => n1740, c => n1741, outb => n1738);
   U2359 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_2_2_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_7_2_port, d => 
                           n370, outb => n1741);
   U2360 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_1_2_port, b
                           => n507, outb => n1740);
   U2361 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_6_2_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_0_2_port, d => 
                           n509, outb => n1739);
   U2362 : aoi22 port map( a => n523, b => n1491, c => n525, d => n1499, outb 
                           => n1737);
   U2363 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_4_2_port, 
                           outb => n1499);
   U2364 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_5_2_port, 
                           outb => n1491);
   U2365 : nand2 port map( a => n527, b => n1507, outb => n1736);
   U2366 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_3_2_port, 
                           outb => n1507);
   U2367 : nand4 port map( a => n1742, b => n1743, c => n1744, d => n1745, outb
                           => load_n_store_RGB_Array_0_n639);
   U2368 : aoi22 port map( a => n1746, b => n1747, c => load_n_store_we_i, d =>
                           load_n_store_lazy_in_0_1_port, outb => n1745);
   U2369 : nor3 port map( a => n1748, b => n1749, c => n1750, outb => n1747);
   U2370 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_26_1_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_31_1_port, d =>
                           n370, outb => n1750);
   U2371 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_25_1_port, 
                           b => n507, outb => n1749);
   U2372 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_30_1_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_24_1_port, d =>
                           n509, outb => n1748);
   U2373 : nor3 port map( a => n1751, b => n1752, c => n512, outb => n1746);
   U2374 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_27_1_port, 
                           b => n513, outb => n1752);
   U2375 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_28_1_port,
                           b => n514, c => 
                           load_n_store_RGB_Array_0_block_ram_r_29_1_port, d =>
                           n515, outb => n1751);
   U2376 : nand4 port map( a => n516, b => n1753, c => n1754, d => n1755, outb 
                           => n1744);
   U2377 : nor3 port map( a => n1756, b => n1757, c => n1758, outb => n1755);
   U2378 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_18_1_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_23_1_port, d =>
                           n370, outb => n1758);
   U2379 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_17_1_port, 
                           b => n507, outb => n1757);
   U2380 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_22_1_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_16_1_port, d =>
                           n509, outb => n1756);
   U2381 : aoi22 port map( a => n523, b => n1759, c => n525, d => n1760, outb 
                           => n1754);
   U2382 : nand2 port map( a => n527, b => n1761, outb => n1753);
   U2383 : nand4 port map( a => n529, b => n1762, c => n1763, d => n1764, outb 
                           => n1743);
   U2384 : nor3 port map( a => n1765, b => n1766, c => n1767, outb => n1764);
   U2385 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_10_1_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_15_1_port, d =>
                           n370, outb => n1767);
   U2386 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_9_1_port, b
                           => n507, outb => n1766);
   U2387 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_14_1_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_8_1_port, d => 
                           n509, outb => n1765);
   U2388 : aoi22 port map( a => n523, b => n1768, c => n525, d => n1769, outb 
                           => n1763);
   U2389 : nand2 port map( a => n527, b => n1437, outb => n1762);
   U2390 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_11_1_port,
                           outb => n1437);
   U2391 : nand4 port map( a => n539, b => n1770, c => n1771, d => n1772, outb 
                           => n1742);
   U2392 : nor3 port map( a => n1773, b => n1774, c => n1775, outb => n1772);
   U2393 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_2_1_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_7_1_port, d => 
                           n370, outb => n1775);
   U2394 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_1_1_port, b
                           => n507, outb => n1774);
   U2395 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_6_1_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_0_1_port, d => 
                           n509, outb => n1773);
   U2396 : aoi22 port map( a => n523, b => n1492, c => n525, d => n1500, outb 
                           => n1771);
   U2397 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_4_1_port, 
                           outb => n1500);
   U2398 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_5_1_port, 
                           outb => n1492);
   U2399 : nand2 port map( a => n527, b => n1508, outb => n1770);
   U2400 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_3_1_port, 
                           outb => n1508);
   U2401 : nand4 port map( a => n1776, b => n1777, c => n1778, d => n1779, outb
                           => load_n_store_RGB_Array_0_n636);
   U2402 : aoi22 port map( a => n1780, b => n1781, c => load_n_store_we_i, d =>
                           load_n_store_lazy_in_0_0_port, outb => n1779);
   U2403 : nor3 port map( a => n1782, b => n1783, c => n1784, outb => n1781);
   U2404 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_26_0_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_31_0_port, d =>
                           n370, outb => n1784);
   U2405 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_25_0_port, 
                           b => n507, outb => n1783);
   U2406 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_30_0_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_24_0_port, d =>
                           n509, outb => n1782);
   U2407 : nor3 port map( a => n1785, b => n1786, c => n512, outb => n1780);
   U2408 : inv port map( inb => n1787, outb => n512);
   U2409 : nor2 port map( a => n371, b => load_n_store_we_i, outb => n1787);
   U2410 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_27_0_port, 
                           b => n513, outb => n1786);
   U2411 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_28_0_port,
                           b => n514, c => 
                           load_n_store_RGB_Array_0_block_ram_r_29_0_port, d =>
                           n515, outb => n1785);
   U2412 : nand4 port map( a => n516, b => n1788, c => n1789, d => n1790, outb 
                           => n1778);
   U2413 : nor3 port map( a => n1791, b => n1792, c => n1793, outb => n1790);
   U2414 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_18_0_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_23_0_port, d =>
                           n370, outb => n1793);
   U2415 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_17_0_port, 
                           b => n507, outb => n1792);
   U2416 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_22_0_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_16_0_port, d =>
                           n509, outb => n1791);
   U2417 : aoi22 port map( a => n523, b => n1794, c => n525, d => n1795, outb 
                           => n1789);
   U2418 : nand2 port map( a => n527, b => n1796, outb => n1788);
   U2419 : nor3 port map( a => load_n_store_s_addr_3_port, b => 
                           load_n_store_we_i, c => n312, outb => n516);
   U2420 : nand4 port map( a => n529, b => n1797, c => n1798, d => n1799, outb 
                           => n1777);
   U2421 : nor3 port map( a => n1800, b => n1801, c => n1802, outb => n1799);
   U2422 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_10_0_port,
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_15_0_port, d =>
                           n370, outb => n1802);
   U2423 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_9_0_port, b
                           => n507, outb => n1801);
   U2424 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_14_0_port,
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_8_0_port, d => 
                           n509, outb => n1800);
   U2425 : aoi22 port map( a => n523, b => n1803, c => n525, d => n1804, outb 
                           => n1798);
   U2426 : nand2 port map( a => n527, b => n1438, outb => n1797);
   U2427 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_11_0_port,
                           outb => n1438);
   U2428 : nor3 port map( a => load_n_store_s_addr_4_port, b => 
                           load_n_store_we_i, c => n315, outb => n529);
   U2429 : nand4 port map( a => n539, b => n1805, c => n1806, d => n1807, outb 
                           => n1776);
   U2430 : nor3 port map( a => n1808, b => n1809, c => n1810, outb => n1807);
   U2431 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_2_0_port, 
                           b => n506, c => 
                           load_n_store_RGB_Array_0_block_ram_r_7_0_port, d => 
                           n370, outb => n1810);
   U2432 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_1_0_port, b
                           => n507, outb => n1809);
   U2433 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_6_0_port, 
                           b => n508, c => 
                           load_n_store_RGB_Array_0_block_ram_r_0_0_port, d => 
                           n509, outb => n1808);
   U2434 : aoi22 port map( a => n523, b => n1493, c => n525, d => n1501, outb 
                           => n1806);
   U2435 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_4_0_port, 
                           outb => n1501);
   U2436 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_5_0_port, 
                           outb => n1493);
   U2437 : nand2 port map( a => n527, b => n1509, outb => n1805);
   U2438 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_3_0_port, 
                           outb => n1509);
   U2439 : nor3 port map( a => load_n_store_s_addr_4_port, b => 
                           load_n_store_we_i, c => load_n_store_s_addr_3_port, 
                           outb => n539);
   U2440 : oai22 port map( a => n215, b => n786, c => n787, d => n1811, outb =>
                           load_n_store_RGB_Array_0_n1162);
   U2441 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_31_7_port,
                           outb => n1811);
   U2442 : oai22 port map( a => n213, b => n786, c => n787, d => n1812, outb =>
                           load_n_store_RGB_Array_0_n1161);
   U2443 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_31_6_port,
                           outb => n1812);
   U2444 : oai22 port map( a => n211, b => n786, c => n787, d => n1813, outb =>
                           load_n_store_RGB_Array_0_n1160);
   U2445 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_31_5_port,
                           outb => n1813);
   U2446 : oai22 port map( a => n209, b => n786, c => n787, d => n1814, outb =>
                           load_n_store_RGB_Array_0_n1159);
   U2447 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_31_4_port,
                           outb => n1814);
   U2448 : oai22 port map( a => n207, b => n786, c => n787, d => n1815, outb =>
                           load_n_store_RGB_Array_0_n1158);
   U2449 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_31_3_port,
                           outb => n1815);
   U2450 : oai22 port map( a => n205, b => n786, c => n787, d => n1816, outb =>
                           load_n_store_RGB_Array_0_n1157);
   U2451 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_31_2_port,
                           outb => n1816);
   U2452 : oai22 port map( a => n203, b => n786, c => n787, d => n1817, outb =>
                           load_n_store_RGB_Array_0_n1156);
   U2453 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_31_1_port,
                           outb => n1817);
   U2454 : oai22 port map( a => n201, b => n786, c => n787, d => n1818, outb =>
                           load_n_store_RGB_Array_0_n1155);
   U2455 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_31_0_port,
                           outb => n1818);
   U2456 : inv port map( inb => n786, outb => n787);
   U2457 : nand2 port map( a => n1819, b => n1476, outb => n786);
   U2458 : oai22 port map( a => n215, b => n796, c => n797, d => n1820, outb =>
                           load_n_store_RGB_Array_0_n1154);
   U2459 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_30_7_port,
                           outb => n1820);
   U2460 : oai22 port map( a => n213, b => n796, c => n797, d => n1821, outb =>
                           load_n_store_RGB_Array_0_n1153);
   U2461 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_30_6_port,
                           outb => n1821);
   U2462 : oai22 port map( a => n211, b => n796, c => n797, d => n1822, outb =>
                           load_n_store_RGB_Array_0_n1152);
   U2463 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_30_5_port,
                           outb => n1822);
   U2464 : oai22 port map( a => n209, b => n796, c => n797, d => n1823, outb =>
                           load_n_store_RGB_Array_0_n1151);
   U2465 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_30_4_port,
                           outb => n1823);
   U2466 : oai22 port map( a => n207, b => n796, c => n797, d => n1824, outb =>
                           load_n_store_RGB_Array_0_n1150);
   U2467 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_30_3_port,
                           outb => n1824);
   U2468 : oai22 port map( a => n205, b => n796, c => n797, d => n1825, outb =>
                           load_n_store_RGB_Array_0_n1149);
   U2469 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_30_2_port,
                           outb => n1825);
   U2470 : oai22 port map( a => n203, b => n796, c => n797, d => n1826, outb =>
                           load_n_store_RGB_Array_0_n1148);
   U2471 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_30_1_port,
                           outb => n1826);
   U2472 : oai22 port map( a => n201, b => n796, c => n797, d => n1827, outb =>
                           load_n_store_RGB_Array_0_n1147);
   U2473 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_30_0_port,
                           outb => n1827);
   U2474 : inv port map( inb => n796, outb => n797);
   U2475 : nand2 port map( a => n1819, b => n1485, outb => n796);
   U2476 : oai22 port map( a => n215, b => n806, c => n807, d => n1828, outb =>
                           load_n_store_RGB_Array_0_n1146);
   U2477 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_29_7_port,
                           outb => n1828);
   U2478 : oai22 port map( a => n213, b => n806, c => n807, d => n1829, outb =>
                           load_n_store_RGB_Array_0_n1145);
   U2479 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_29_6_port,
                           outb => n1829);
   U2480 : oai22 port map( a => n211, b => n806, c => n807, d => n1830, outb =>
                           load_n_store_RGB_Array_0_n1144);
   U2481 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_29_5_port,
                           outb => n1830);
   U2482 : oai22 port map( a => n209, b => n806, c => n807, d => n1831, outb =>
                           load_n_store_RGB_Array_0_n1143);
   U2483 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_29_4_port,
                           outb => n1831);
   U2484 : oai22 port map( a => n207, b => n806, c => n807, d => n1832, outb =>
                           load_n_store_RGB_Array_0_n1142);
   U2485 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_29_3_port,
                           outb => n1832);
   U2486 : oai22 port map( a => n205, b => n806, c => n807, d => n1833, outb =>
                           load_n_store_RGB_Array_0_n1141);
   U2487 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_29_2_port,
                           outb => n1833);
   U2488 : oai22 port map( a => n203, b => n806, c => n807, d => n1834, outb =>
                           load_n_store_RGB_Array_0_n1140);
   U2489 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_29_1_port,
                           outb => n1834);
   U2490 : oai22 port map( a => n201, b => n806, c => n807, d => n1835, outb =>
                           load_n_store_RGB_Array_0_n1139);
   U2491 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_29_0_port,
                           outb => n1835);
   U2492 : inv port map( inb => n806, outb => n807);
   U2493 : nand2 port map( a => n1819, b => n523, outb => n806);
   U2494 : oai22 port map( a => n215, b => n816, c => n817, d => n1836, outb =>
                           load_n_store_RGB_Array_0_n1138);
   U2495 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_28_7_port,
                           outb => n1836);
   U2496 : oai22 port map( a => n213, b => n816, c => n817, d => n1837, outb =>
                           load_n_store_RGB_Array_0_n1137);
   U2497 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_28_6_port,
                           outb => n1837);
   U2498 : oai22 port map( a => n211, b => n816, c => n817, d => n1838, outb =>
                           load_n_store_RGB_Array_0_n1136);
   U2499 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_28_5_port,
                           outb => n1838);
   U2500 : oai22 port map( a => n209, b => n816, c => n817, d => n1839, outb =>
                           load_n_store_RGB_Array_0_n1135);
   U2501 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_28_4_port,
                           outb => n1839);
   U2502 : oai22 port map( a => n207, b => n816, c => n817, d => n1840, outb =>
                           load_n_store_RGB_Array_0_n1134);
   U2503 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_28_3_port,
                           outb => n1840);
   U2504 : oai22 port map( a => n205, b => n816, c => n817, d => n1841, outb =>
                           load_n_store_RGB_Array_0_n1133);
   U2505 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_28_2_port,
                           outb => n1841);
   U2506 : oai22 port map( a => n203, b => n816, c => n817, d => n1842, outb =>
                           load_n_store_RGB_Array_0_n1132);
   U2507 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_28_1_port,
                           outb => n1842);
   U2508 : oai22 port map( a => n201, b => n816, c => n817, d => n1843, outb =>
                           load_n_store_RGB_Array_0_n1131);
   U2509 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_28_0_port,
                           outb => n1843);
   U2510 : inv port map( inb => n816, outb => n817);
   U2511 : nand2 port map( a => n1819, b => n525, outb => n816);
   U2512 : oai22 port map( a => n215, b => n826, c => n827, d => n1844, outb =>
                           load_n_store_RGB_Array_0_n1130);
   U2513 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_27_7_port,
                           outb => n1844);
   U2514 : oai22 port map( a => n213, b => n826, c => n827, d => n1845, outb =>
                           load_n_store_RGB_Array_0_n1129);
   U2515 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_27_6_port,
                           outb => n1845);
   U2516 : oai22 port map( a => n211, b => n826, c => n827, d => n1846, outb =>
                           load_n_store_RGB_Array_0_n1128);
   U2517 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_27_5_port,
                           outb => n1846);
   U2518 : oai22 port map( a => n209, b => n826, c => n827, d => n1847, outb =>
                           load_n_store_RGB_Array_0_n1127);
   U2519 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_27_4_port,
                           outb => n1847);
   U2520 : oai22 port map( a => n207, b => n826, c => n827, d => n1848, outb =>
                           load_n_store_RGB_Array_0_n1126);
   U2521 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_27_3_port,
                           outb => n1848);
   U2522 : oai22 port map( a => n205, b => n826, c => n827, d => n1849, outb =>
                           load_n_store_RGB_Array_0_n1125);
   U2523 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_27_2_port,
                           outb => n1849);
   U2524 : oai22 port map( a => n203, b => n826, c => n827, d => n1850, outb =>
                           load_n_store_RGB_Array_0_n1124);
   U2525 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_27_1_port,
                           outb => n1850);
   U2526 : oai22 port map( a => n201, b => n826, c => n827, d => n1851, outb =>
                           load_n_store_RGB_Array_0_n1123);
   U2527 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_27_0_port,
                           outb => n1851);
   U2528 : inv port map( inb => n826, outb => n827);
   U2529 : nand2 port map( a => n1819, b => n527, outb => n826);
   U2530 : oai22 port map( a => n215, b => n836, c => n837, d => n1852, outb =>
                           load_n_store_RGB_Array_0_n1122);
   U2531 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_26_7_port,
                           outb => n1852);
   U2532 : oai22 port map( a => n213, b => n836, c => n837, d => n1853, outb =>
                           load_n_store_RGB_Array_0_n1121);
   U2533 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_26_6_port,
                           outb => n1853);
   U2534 : oai22 port map( a => n211, b => n836, c => n837, d => n1854, outb =>
                           load_n_store_RGB_Array_0_n1120);
   U2535 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_26_5_port,
                           outb => n1854);
   U2536 : oai22 port map( a => n209, b => n836, c => n837, d => n1855, outb =>
                           load_n_store_RGB_Array_0_n1119);
   U2537 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_26_4_port,
                           outb => n1855);
   U2538 : oai22 port map( a => n207, b => n836, c => n837, d => n1856, outb =>
                           load_n_store_RGB_Array_0_n1118);
   U2539 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_26_3_port,
                           outb => n1856);
   U2540 : oai22 port map( a => n205, b => n836, c => n837, d => n1857, outb =>
                           load_n_store_RGB_Array_0_n1117);
   U2541 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_26_2_port,
                           outb => n1857);
   U2542 : oai22 port map( a => n203, b => n836, c => n837, d => n1858, outb =>
                           load_n_store_RGB_Array_0_n1116);
   U2543 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_26_1_port,
                           outb => n1858);
   U2544 : oai22 port map( a => n201, b => n836, c => n837, d => n1859, outb =>
                           load_n_store_RGB_Array_0_n1115);
   U2545 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_26_0_port,
                           outb => n1859);
   U2546 : inv port map( inb => n836, outb => n837);
   U2547 : nand2 port map( a => n1819, b => n1447, outb => n836);
   U2548 : oai22 port map( a => n215, b => n846, c => n847, d => n1860, outb =>
                           load_n_store_RGB_Array_0_n1114);
   U2549 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_25_7_port,
                           outb => n1860);
   U2550 : oai22 port map( a => n213, b => n846, c => n847, d => n1861, outb =>
                           load_n_store_RGB_Array_0_n1113);
   U2551 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_25_6_port,
                           outb => n1861);
   U2552 : oai22 port map( a => n211, b => n846, c => n847, d => n1862, outb =>
                           load_n_store_RGB_Array_0_n1112);
   U2553 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_25_5_port,
                           outb => n1862);
   U2554 : oai22 port map( a => n209, b => n846, c => n847, d => n1863, outb =>
                           load_n_store_RGB_Array_0_n1111);
   U2555 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_25_4_port,
                           outb => n1863);
   U2556 : oai22 port map( a => n207, b => n846, c => n847, d => n1864, outb =>
                           load_n_store_RGB_Array_0_n1110);
   U2557 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_25_3_port,
                           outb => n1864);
   U2558 : oai22 port map( a => n205, b => n846, c => n847, d => n1865, outb =>
                           load_n_store_RGB_Array_0_n1109);
   U2559 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_25_2_port,
                           outb => n1865);
   U2560 : oai22 port map( a => n203, b => n846, c => n847, d => n1866, outb =>
                           load_n_store_RGB_Array_0_n1108);
   U2561 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_25_1_port,
                           outb => n1866);
   U2562 : oai22 port map( a => n201, b => n846, c => n847, d => n1867, outb =>
                           load_n_store_RGB_Array_0_n1107);
   U2563 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_25_0_port,
                           outb => n1867);
   U2564 : inv port map( inb => n846, outb => n847);
   U2565 : nand2 port map( a => n1819, b => n1457, outb => n846);
   U2566 : oai22 port map( a => n215, b => n856, c => n857, d => n1868, outb =>
                           load_n_store_RGB_Array_0_n1106);
   U2567 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_24_7_port,
                           outb => n1868);
   U2568 : oai22 port map( a => n213, b => n856, c => n857, d => n1869, outb =>
                           load_n_store_RGB_Array_0_n1105);
   U2569 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_24_6_port,
                           outb => n1869);
   U2570 : oai22 port map( a => n211, b => n856, c => n857, d => n1870, outb =>
                           load_n_store_RGB_Array_0_n1104);
   U2571 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_24_5_port,
                           outb => n1870);
   U2572 : oai22 port map( a => n209, b => n856, c => n857, d => n1871, outb =>
                           load_n_store_RGB_Array_0_n1103);
   U2573 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_24_4_port,
                           outb => n1871);
   U2574 : oai22 port map( a => n207, b => n856, c => n857, d => n1872, outb =>
                           load_n_store_RGB_Array_0_n1102);
   U2575 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_24_3_port,
                           outb => n1872);
   U2576 : oai22 port map( a => n205, b => n856, c => n857, d => n1873, outb =>
                           load_n_store_RGB_Array_0_n1101);
   U2577 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_24_2_port,
                           outb => n1873);
   U2578 : oai22 port map( a => n203, b => n856, c => n857, d => n1874, outb =>
                           load_n_store_RGB_Array_0_n1100);
   U2579 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_24_1_port,
                           outb => n1874);
   U2580 : oai22 port map( a => n201, b => n856, c => n857, d => n1875, outb =>
                           load_n_store_RGB_Array_0_n1099);
   U2581 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_24_0_port,
                           outb => n1875);
   U2582 : inv port map( inb => n856, outb => n857);
   U2583 : nand2 port map( a => n1819, b => n1466, outb => n856);
   U2584 : nor2 port map( a => n1534, b => n371, outb => n1819);
   U2585 : nand2 port map( a => load_n_store_s_addr_4_port, b => 
                           load_n_store_s_addr_3_port, outb => n371);
   U2586 : oai22 port map( a => n215, b => n866, c => n867, d => n1876, outb =>
                           load_n_store_RGB_Array_0_n1098);
   U2587 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_23_7_port,
                           outb => n1876);
   U2588 : oai22 port map( a => n213, b => n866, c => n867, d => n1877, outb =>
                           load_n_store_RGB_Array_0_n1097);
   U2589 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_23_6_port,
                           outb => n1877);
   U2590 : oai22 port map( a => n211, b => n866, c => n867, d => n1878, outb =>
                           load_n_store_RGB_Array_0_n1096);
   U2591 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_23_5_port,
                           outb => n1878);
   U2592 : oai22 port map( a => n209, b => n866, c => n867, d => n1879, outb =>
                           load_n_store_RGB_Array_0_n1095);
   U2593 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_23_4_port,
                           outb => n1879);
   U2594 : oai22 port map( a => n207, b => n866, c => n867, d => n1880, outb =>
                           load_n_store_RGB_Array_0_n1094);
   U2595 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_23_3_port,
                           outb => n1880);
   U2596 : oai22 port map( a => n205, b => n866, c => n867, d => n1881, outb =>
                           load_n_store_RGB_Array_0_n1093);
   U2597 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_23_2_port,
                           outb => n1881);
   U2598 : oai22 port map( a => n203, b => n866, c => n867, d => n1882, outb =>
                           load_n_store_RGB_Array_0_n1092);
   U2599 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_23_1_port,
                           outb => n1882);
   U2600 : oai22 port map( a => n201, b => n866, c => n867, d => n1883, outb =>
                           load_n_store_RGB_Array_0_n1091);
   U2601 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_23_0_port,
                           outb => n1883);
   U2602 : inv port map( inb => n866, outb => n867);
   U2603 : nand2 port map( a => n1884, b => n1476, outb => n866);
   U2604 : oai22 port map( a => n215, b => n876, c => n877, d => n1885, outb =>
                           load_n_store_RGB_Array_0_n1090);
   U2605 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_22_7_port,
                           outb => n1885);
   U2606 : oai22 port map( a => n213, b => n876, c => n877, d => n1886, outb =>
                           load_n_store_RGB_Array_0_n1089);
   U2607 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_22_6_port,
                           outb => n1886);
   U2608 : oai22 port map( a => n211, b => n876, c => n877, d => n1887, outb =>
                           load_n_store_RGB_Array_0_n1088);
   U2609 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_22_5_port,
                           outb => n1887);
   U2610 : oai22 port map( a => n209, b => n876, c => n877, d => n1888, outb =>
                           load_n_store_RGB_Array_0_n1087);
   U2611 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_22_4_port,
                           outb => n1888);
   U2612 : oai22 port map( a => n207, b => n876, c => n877, d => n1889, outb =>
                           load_n_store_RGB_Array_0_n1086);
   U2613 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_22_3_port,
                           outb => n1889);
   U2614 : oai22 port map( a => n205, b => n876, c => n877, d => n1890, outb =>
                           load_n_store_RGB_Array_0_n1085);
   U2615 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_22_2_port,
                           outb => n1890);
   U2616 : oai22 port map( a => n203, b => n876, c => n877, d => n1891, outb =>
                           load_n_store_RGB_Array_0_n1084);
   U2617 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_22_1_port,
                           outb => n1891);
   U2618 : oai22 port map( a => n201, b => n876, c => n877, d => n1892, outb =>
                           load_n_store_RGB_Array_0_n1083);
   U2619 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_22_0_port,
                           outb => n1892);
   U2620 : inv port map( inb => n876, outb => n877);
   U2621 : nand2 port map( a => n1884, b => n1485, outb => n876);
   U2622 : oai22 port map( a => n215, b => n886, c => n887, d => n1552, outb =>
                           load_n_store_RGB_Array_0_n1082);
   U2623 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_21_7_port,
                           outb => n1552);
   U2624 : oai22 port map( a => n213, b => n886, c => n887, d => n1587, outb =>
                           load_n_store_RGB_Array_0_n1081);
   U2625 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_21_6_port,
                           outb => n1587);
   U2626 : oai22 port map( a => n211, b => n886, c => n887, d => n1622, outb =>
                           load_n_store_RGB_Array_0_n1080);
   U2627 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_21_5_port,
                           outb => n1622);
   U2628 : oai22 port map( a => n209, b => n886, c => n887, d => n1657, outb =>
                           load_n_store_RGB_Array_0_n1079);
   U2629 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_21_4_port,
                           outb => n1657);
   U2630 : oai22 port map( a => n207, b => n886, c => n887, d => n1691, outb =>
                           load_n_store_RGB_Array_0_n1078);
   U2631 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_21_3_port,
                           outb => n1691);
   U2632 : oai22 port map( a => n205, b => n886, c => n887, d => n1725, outb =>
                           load_n_store_RGB_Array_0_n1077);
   U2633 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_21_2_port,
                           outb => n1725);
   U2634 : oai22 port map( a => n203, b => n886, c => n887, d => n1759, outb =>
                           load_n_store_RGB_Array_0_n1076);
   U2635 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_21_1_port,
                           outb => n1759);
   U2636 : oai22 port map( a => n201, b => n886, c => n887, d => n1794, outb =>
                           load_n_store_RGB_Array_0_n1075);
   U2637 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_21_0_port,
                           outb => n1794);
   U2638 : inv port map( inb => n886, outb => n887);
   U2639 : nand2 port map( a => n1884, b => n523, outb => n886);
   U2640 : oai22 port map( a => n215, b => n888, c => n889, d => n1553, outb =>
                           load_n_store_RGB_Array_0_n1074);
   U2641 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_20_7_port,
                           outb => n1553);
   U2642 : oai22 port map( a => n213, b => n888, c => n889, d => n1588, outb =>
                           load_n_store_RGB_Array_0_n1073);
   U2643 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_20_6_port,
                           outb => n1588);
   U2644 : oai22 port map( a => n211, b => n888, c => n889, d => n1623, outb =>
                           load_n_store_RGB_Array_0_n1072);
   U2645 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_20_5_port,
                           outb => n1623);
   U2646 : oai22 port map( a => n209, b => n888, c => n889, d => n1658, outb =>
                           load_n_store_RGB_Array_0_n1071);
   U2647 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_20_4_port,
                           outb => n1658);
   U2648 : oai22 port map( a => n207, b => n888, c => n889, d => n1692, outb =>
                           load_n_store_RGB_Array_0_n1070);
   U2649 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_20_3_port,
                           outb => n1692);
   U2650 : oai22 port map( a => n205, b => n888, c => n889, d => n1726, outb =>
                           load_n_store_RGB_Array_0_n1069);
   U2651 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_20_2_port,
                           outb => n1726);
   U2652 : oai22 port map( a => n203, b => n888, c => n889, d => n1760, outb =>
                           load_n_store_RGB_Array_0_n1068);
   U2653 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_20_1_port,
                           outb => n1760);
   U2654 : oai22 port map( a => n201, b => n888, c => n889, d => n1795, outb =>
                           load_n_store_RGB_Array_0_n1067);
   U2655 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_20_0_port,
                           outb => n1795);
   U2656 : inv port map( inb => n888, outb => n889);
   U2657 : nand2 port map( a => n1884, b => n525, outb => n888);
   U2658 : oai22 port map( a => n215, b => n890, c => n891, d => n1554, outb =>
                           load_n_store_RGB_Array_0_n1066);
   U2659 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_19_7_port,
                           outb => n1554);
   U2660 : oai22 port map( a => n213, b => n890, c => n891, d => n1589, outb =>
                           load_n_store_RGB_Array_0_n1065);
   U2661 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_19_6_port,
                           outb => n1589);
   U2662 : oai22 port map( a => n211, b => n890, c => n891, d => n1624, outb =>
                           load_n_store_RGB_Array_0_n1064);
   U2663 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_19_5_port,
                           outb => n1624);
   U2664 : oai22 port map( a => n209, b => n890, c => n891, d => n1659, outb =>
                           load_n_store_RGB_Array_0_n1063);
   U2665 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_19_4_port,
                           outb => n1659);
   U2666 : oai22 port map( a => n207, b => n890, c => n891, d => n1693, outb =>
                           load_n_store_RGB_Array_0_n1062);
   U2667 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_19_3_port,
                           outb => n1693);
   U2668 : oai22 port map( a => n205, b => n890, c => n891, d => n1727, outb =>
                           load_n_store_RGB_Array_0_n1061);
   U2669 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_19_2_port,
                           outb => n1727);
   U2670 : oai22 port map( a => n203, b => n890, c => n891, d => n1761, outb =>
                           load_n_store_RGB_Array_0_n1060);
   U2671 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_19_1_port,
                           outb => n1761);
   U2672 : oai22 port map( a => n201, b => n890, c => n891, d => n1796, outb =>
                           load_n_store_RGB_Array_0_n1059);
   U2673 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_19_0_port,
                           outb => n1796);
   U2674 : inv port map( inb => n890, outb => n891);
   U2675 : nand2 port map( a => n1884, b => n527, outb => n890);
   U2676 : oai22 port map( a => n215, b => n892, c => n893, d => n1893, outb =>
                           load_n_store_RGB_Array_0_n1058);
   U2677 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_18_7_port,
                           outb => n1893);
   U2678 : oai22 port map( a => n213, b => n892, c => n893, d => n1894, outb =>
                           load_n_store_RGB_Array_0_n1057);
   U2679 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_18_6_port,
                           outb => n1894);
   U2680 : oai22 port map( a => n211, b => n892, c => n893, d => n1895, outb =>
                           load_n_store_RGB_Array_0_n1056);
   U2681 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_18_5_port,
                           outb => n1895);
   U2682 : oai22 port map( a => n209, b => n892, c => n893, d => n1896, outb =>
                           load_n_store_RGB_Array_0_n1055);
   U2683 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_18_4_port,
                           outb => n1896);
   U2684 : oai22 port map( a => n207, b => n892, c => n893, d => n1897, outb =>
                           load_n_store_RGB_Array_0_n1054);
   U2685 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_18_3_port,
                           outb => n1897);
   U2686 : oai22 port map( a => n205, b => n892, c => n893, d => n1898, outb =>
                           load_n_store_RGB_Array_0_n1053);
   U2687 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_18_2_port,
                           outb => n1898);
   U2688 : oai22 port map( a => n203, b => n892, c => n893, d => n1899, outb =>
                           load_n_store_RGB_Array_0_n1052);
   U2689 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_18_1_port,
                           outb => n1899);
   U2690 : oai22 port map( a => n201, b => n892, c => n893, d => n1900, outb =>
                           load_n_store_RGB_Array_0_n1051);
   U2691 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_18_0_port,
                           outb => n1900);
   U2692 : inv port map( inb => n892, outb => n893);
   U2693 : nand2 port map( a => n1884, b => n1447, outb => n892);
   U2694 : inv port map( inb => n506, outb => n1447);
   U2695 : nand3 port map( a => n304, b => n363, c => 
                           load_n_store_s_addr_1_port, outb => n506);
   U2696 : oai22 port map( a => n215, b => n902, c => n903, d => n1901, outb =>
                           load_n_store_RGB_Array_0_n1050);
   U2697 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_17_7_port,
                           outb => n1901);
   U2698 : oai22 port map( a => n213, b => n902, c => n903, d => n1902, outb =>
                           load_n_store_RGB_Array_0_n1049);
   U2699 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_17_6_port,
                           outb => n1902);
   U2700 : oai22 port map( a => n211, b => n902, c => n903, d => n1903, outb =>
                           load_n_store_RGB_Array_0_n1048);
   U2701 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_17_5_port,
                           outb => n1903);
   U2702 : oai22 port map( a => n209, b => n902, c => n903, d => n1904, outb =>
                           load_n_store_RGB_Array_0_n1047);
   U2703 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_17_4_port,
                           outb => n1904);
   U2704 : oai22 port map( a => n207, b => n902, c => n903, d => n1905, outb =>
                           load_n_store_RGB_Array_0_n1046);
   U2705 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_17_3_port,
                           outb => n1905);
   U2706 : oai22 port map( a => n205, b => n902, c => n903, d => n1906, outb =>
                           load_n_store_RGB_Array_0_n1045);
   U2707 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_17_2_port,
                           outb => n1906);
   U2708 : oai22 port map( a => n203, b => n902, c => n903, d => n1907, outb =>
                           load_n_store_RGB_Array_0_n1044);
   U2709 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_17_1_port,
                           outb => n1907);
   U2710 : oai22 port map( a => n201, b => n902, c => n903, d => n1908, outb =>
                           load_n_store_RGB_Array_0_n1043);
   U2711 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_17_0_port,
                           outb => n1908);
   U2712 : inv port map( inb => n902, outb => n903);
   U2713 : nand2 port map( a => n1884, b => n1457, outb => n902);
   U2714 : inv port map( inb => n507, outb => n1457);
   U2715 : nand3 port map( a => n359, b => n363, c => 
                           load_n_store_s_addr_0_port, outb => n507);
   U2716 : oai22 port map( a => n215, b => n912, c => n913, d => n1909, outb =>
                           load_n_store_RGB_Array_0_n1042);
   U2717 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_16_7_port,
                           outb => n1909);
   U2718 : oai22 port map( a => n213, b => n912, c => n913, d => n1910, outb =>
                           load_n_store_RGB_Array_0_n1041);
   U2719 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_16_6_port,
                           outb => n1910);
   U2720 : oai22 port map( a => n211, b => n912, c => n913, d => n1911, outb =>
                           load_n_store_RGB_Array_0_n1040);
   U2721 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_16_5_port,
                           outb => n1911);
   U2722 : oai22 port map( a => n209, b => n912, c => n913, d => n1912, outb =>
                           load_n_store_RGB_Array_0_n1039);
   U2723 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_16_4_port,
                           outb => n1912);
   U2724 : oai22 port map( a => n207, b => n912, c => n913, d => n1913, outb =>
                           load_n_store_RGB_Array_0_n1038);
   U2725 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_16_3_port,
                           outb => n1913);
   U2726 : oai22 port map( a => n205, b => n912, c => n913, d => n1914, outb =>
                           load_n_store_RGB_Array_0_n1037);
   U2727 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_16_2_port,
                           outb => n1914);
   U2728 : oai22 port map( a => n203, b => n912, c => n913, d => n1915, outb =>
                           load_n_store_RGB_Array_0_n1036);
   U2729 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_16_1_port,
                           outb => n1915);
   U2730 : oai22 port map( a => n201, b => n912, c => n913, d => n1916, outb =>
                           load_n_store_RGB_Array_0_n1035);
   U2731 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_16_0_port,
                           outb => n1916);
   U2732 : inv port map( inb => n912, outb => n913);
   U2733 : nand2 port map( a => n1884, b => n1466, outb => n912);
   U2734 : inv port map( inb => n509, outb => n1466);
   U2735 : nand3 port map( a => n359, b => n363, c => n304, outb => n509);
   U2736 : nor3 port map( a => n312, b => load_n_store_s_addr_3_port, c => 
                           n1534, outb => n1884);
   U2737 : inv port map( inb => load_n_store_s_addr_4_port, outb => n312);
   U2738 : oai22 port map( a => n215, b => n922, c => n923, d => n1917, outb =>
                           load_n_store_RGB_Array_0_n1034);
   U2739 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_15_7_port,
                           outb => n1917);
   U2740 : oai22 port map( a => n213, b => n922, c => n923, d => n1918, outb =>
                           load_n_store_RGB_Array_0_n1033);
   U2741 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_15_6_port,
                           outb => n1918);
   U2742 : oai22 port map( a => n211, b => n922, c => n923, d => n1919, outb =>
                           load_n_store_RGB_Array_0_n1032);
   U2743 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_15_5_port,
                           outb => n1919);
   U2744 : oai22 port map( a => n209, b => n922, c => n923, d => n1920, outb =>
                           load_n_store_RGB_Array_0_n1031);
   U2745 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_15_4_port,
                           outb => n1920);
   U2746 : oai22 port map( a => n207, b => n922, c => n923, d => n1921, outb =>
                           load_n_store_RGB_Array_0_n1030);
   U2747 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_15_3_port,
                           outb => n1921);
   U2748 : oai22 port map( a => n205, b => n922, c => n923, d => n1922, outb =>
                           load_n_store_RGB_Array_0_n1029);
   U2749 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_15_2_port,
                           outb => n1922);
   U2750 : oai22 port map( a => n203, b => n922, c => n923, d => n1923, outb =>
                           load_n_store_RGB_Array_0_n1028);
   U2751 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_15_1_port,
                           outb => n1923);
   U2752 : oai22 port map( a => n201, b => n922, c => n923, d => n1924, outb =>
                           load_n_store_RGB_Array_0_n1027);
   U2753 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_15_0_port,
                           outb => n1924);
   U2754 : inv port map( inb => n922, outb => n923);
   U2755 : nand2 port map( a => n1448, b => n1476, outb => n922);
   U2756 : inv port map( inb => n370, outb => n1476);
   U2757 : nand3 port map( a => load_n_store_s_addr_1_port, b => 
                           load_n_store_s_addr_0_port, c => 
                           load_n_store_s_addr_2_port, outb => n370);
   U2758 : oai22 port map( a => n215, b => n932, c => n933, d => n1925, outb =>
                           load_n_store_RGB_Array_0_n1026);
   U2759 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_14_7_port,
                           outb => n1925);
   U2760 : oai22 port map( a => n213, b => n932, c => n933, d => n1926, outb =>
                           load_n_store_RGB_Array_0_n1025);
   U2761 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_14_6_port,
                           outb => n1926);
   U2762 : oai22 port map( a => n211, b => n932, c => n933, d => n1927, outb =>
                           load_n_store_RGB_Array_0_n1024);
   U2763 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_14_5_port,
                           outb => n1927);
   U2764 : oai22 port map( a => n209, b => n932, c => n933, d => n1928, outb =>
                           load_n_store_RGB_Array_0_n1023);
   U2765 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_14_4_port,
                           outb => n1928);
   U2766 : oai22 port map( a => n207, b => n932, c => n933, d => n1929, outb =>
                           load_n_store_RGB_Array_0_n1022);
   U2767 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_14_3_port,
                           outb => n1929);
   U2768 : oai22 port map( a => n205, b => n932, c => n933, d => n1930, outb =>
                           load_n_store_RGB_Array_0_n1021);
   U2769 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_14_2_port,
                           outb => n1930);
   U2770 : oai22 port map( a => n203, b => n932, c => n933, d => n1931, outb =>
                           load_n_store_RGB_Array_0_n1020);
   U2771 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_14_1_port,
                           outb => n1931);
   U2772 : oai22 port map( a => n201, b => n932, c => n933, d => n1932, outb =>
                           load_n_store_RGB_Array_0_n1019);
   U2773 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_14_0_port,
                           outb => n1932);
   U2774 : inv port map( inb => n932, outb => n933);
   U2775 : nand2 port map( a => n1485, b => n1448, outb => n932);
   U2776 : inv port map( inb => n508, outb => n1485);
   U2777 : nand3 port map( a => load_n_store_s_addr_1_port, b => n304, c => 
                           load_n_store_s_addr_2_port, outb => n508);
   U2778 : oai22 port map( a => n215, b => n942, c => n943, d => n1561, outb =>
                           load_n_store_RGB_Array_0_n1018);
   U2779 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_13_7_port,
                           outb => n1561);
   U2780 : oai22 port map( a => n213, b => n942, c => n943, d => n1596, outb =>
                           load_n_store_RGB_Array_0_n1017);
   U2781 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_13_6_port,
                           outb => n1596);
   U2782 : oai22 port map( a => n211, b => n942, c => n943, d => n1631, outb =>
                           load_n_store_RGB_Array_0_n1016);
   U2783 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_13_5_port,
                           outb => n1631);
   U2784 : oai22 port map( a => n209, b => n942, c => n943, d => n1666, outb =>
                           load_n_store_RGB_Array_0_n1015);
   U2785 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_13_4_port,
                           outb => n1666);
   U2786 : oai22 port map( a => n207, b => n942, c => n943, d => n1700, outb =>
                           load_n_store_RGB_Array_0_n1014);
   U2787 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_13_3_port,
                           outb => n1700);
   U2788 : oai22 port map( a => n205, b => n942, c => n943, d => n1734, outb =>
                           load_n_store_RGB_Array_0_n1013);
   U2789 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_13_2_port,
                           outb => n1734);
   U2790 : oai22 port map( a => n203, b => n942, c => n943, d => n1768, outb =>
                           load_n_store_RGB_Array_0_n1012);
   U2791 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_13_1_port,
                           outb => n1768);
   U2792 : oai22 port map( a => n201, b => n942, c => n943, d => n1803, outb =>
                           load_n_store_RGB_Array_0_n1011);
   U2793 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_13_0_port,
                           outb => n1803);
   U2794 : inv port map( inb => n942, outb => n943);
   U2795 : nand2 port map( a => n523, b => n1448, outb => n942);
   U2796 : inv port map( inb => n515, outb => n523);
   U2797 : nand3 port map( a => load_n_store_s_addr_0_port, b => n359, c => 
                           load_n_store_s_addr_2_port, outb => n515);
   U2798 : oai22 port map( a => n215, b => n944, c => n945, d => n1562, outb =>
                           load_n_store_RGB_Array_0_n1010);
   U2799 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_12_7_port,
                           outb => n1562);
   U2800 : oai22 port map( a => n213, b => n944, c => n945, d => n1597, outb =>
                           load_n_store_RGB_Array_0_n1009);
   U2801 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_12_6_port,
                           outb => n1597);
   U2802 : oai22 port map( a => n211, b => n944, c => n945, d => n1632, outb =>
                           load_n_store_RGB_Array_0_n1008);
   U2803 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_12_5_port,
                           outb => n1632);
   U2804 : oai22 port map( a => n209, b => n944, c => n945, d => n1667, outb =>
                           load_n_store_RGB_Array_0_n1007);
   U2805 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_12_4_port,
                           outb => n1667);
   U2806 : inv port map( inb => load_n_store_lazy_in_0_4_port, outb => n209);
   U2807 : oai22 port map( a => n207, b => n944, c => n945, d => n1701, outb =>
                           load_n_store_RGB_Array_0_n1006);
   U2808 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_12_3_port,
                           outb => n1701);
   U2809 : inv port map( inb => load_n_store_lazy_in_0_3_port, outb => n207);
   U2810 : oai22 port map( a => n205, b => n944, c => n945, d => n1735, outb =>
                           load_n_store_RGB_Array_0_n1005);
   U2811 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_12_2_port,
                           outb => n1735);
   U2812 : inv port map( inb => load_n_store_lazy_in_0_2_port, outb => n205);
   U2813 : oai22 port map( a => n203, b => n944, c => n945, d => n1769, outb =>
                           load_n_store_RGB_Array_0_n1004);
   U2814 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_12_1_port,
                           outb => n1769);
   U2815 : inv port map( inb => load_n_store_lazy_in_0_1_port, outb => n203);
   U2816 : oai22 port map( a => n201, b => n944, c => n945, d => n1804, outb =>
                           load_n_store_RGB_Array_0_n1003);
   U2817 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_12_0_port,
                           outb => n1804);
   U2818 : inv port map( inb => n944, outb => n945);
   U2819 : nand2 port map( a => n525, b => n1448, outb => n944);
   U2820 : inv port map( inb => n514, outb => n525);
   U2821 : nand3 port map( a => n304, b => n359, c => 
                           load_n_store_s_addr_2_port, outb => n514);
   U2822 : inv port map( inb => load_n_store_s_addr_1_port, outb => n359);
   U2823 : inv port map( inb => load_n_store_s_addr_0_port, outb => n304);
   U2824 : inv port map( inb => load_n_store_lazy_in_0_0_port, outb => n201);
   U2825 : oai22 port map( a => n215, b => n380, c => n381, d => n1563, outb =>
                           load_n_store_RGB_Array_0_n1002);
   U2826 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_11_7_port,
                           outb => n1563);
   U2827 : inv port map( inb => load_n_store_lazy_in_0_7_port, outb => n215);
   U2828 : oai22 port map( a => n213, b => n380, c => n381, d => n1598, outb =>
                           load_n_store_RGB_Array_0_n1001);
   U2829 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_11_6_port,
                           outb => n1598);
   U2830 : inv port map( inb => load_n_store_lazy_in_0_6_port, outb => n213);
   U2831 : oai22 port map( a => n211, b => n380, c => n381, d => n1633, outb =>
                           load_n_store_RGB_Array_0_n1000);
   U2832 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_11_5_port,
                           outb => n1633);
   U2833 : inv port map( inb => n380, outb => n381);
   U2834 : nand2 port map( a => n1448, b => n527, outb => n380);
   U2835 : inv port map( inb => n513, outb => n527);
   U2836 : nand3 port map( a => load_n_store_s_addr_0_port, b => n363, c => 
                           load_n_store_s_addr_1_port, outb => n513);
   U2837 : inv port map( inb => load_n_store_s_addr_2_port, outb => n363);
   U2838 : nor3 port map( a => n315, b => load_n_store_s_addr_4_port, c => 
                           n1534, outb => n1448);
   U2839 : inv port map( inb => load_n_store_we_i, outb => n1534);
   U2840 : inv port map( inb => load_n_store_s_addr_3_port, outb => n315);
   U2841 : inv port map( inb => load_n_store_lazy_in_0_5_port, outb => n211);
   U2842 : nand4 port map( a => n1933, b => n1934, c => n1935, d => n1936, outb
                           => display_out_n535);
   U2843 : nor3 port map( a => n1937, b => n1938, c => n1939, outb => n1936);
   U2844 : nand2 port map( a => n1940, b => display_out_hub_out_sm_0_port, outb
                           => n1935);
   U2845 : nand3 port map( a => n1941, b => n1942, c => n1943, outb => n1933);
   U2846 : oai22 port map( a => n1940, b => n1944, c => n1945, d => n1946, outb
                           => display_out_n534);
   U2847 : nor2 port map( a => n1947, b => n1948, outb => n1944);
   U2848 : nor3 port map( a => n1949, b => reg_hub_f, c => n1950, outb => n1948
                           );
   U2849 : inv port map( inb => mem_hub_f, outb => n1950);
   U2850 : oai22 port map( a => n1951, b => n1952, c => n1953, d => n1954, outb
                           => display_out_n533);
   U2851 : inv port map( inb => display_out_h_col_1_port, outb => n1953);
   U2852 : oai22 port map( a => n1955, b => n1956, c => n1957, d => n1958, outb
                           => display_out_n532);
   U2853 : nor2 port map( a => n1959, b => n1960, outb => n1957);
   U2854 : inv port map( inb => n1961, outb => n1960);
   U2855 : nand4 port map( a => n1962, b => n1963, c => n1964, d => n1934, outb
                           => display_out_n531);
   U2856 : inv port map( inb => n1965, outb => n1934);
   U2857 : nand2 port map( a => n1940, b => display_out_hub_out_sm_1_port, outb
                           => n1964);
   U2858 : inv port map( inb => n1946, outb => n1940);
   U2859 : nand3 port map( a => n1966, b => n1967, c => n1968, outb => n1946);
   U2860 : nand2 port map( a => n1941, b => n1969, outb => n1963);
   U2861 : oai22 port map( a => n235, b => n1970, c => n1971, d => n1972, outb 
                           => display_out_n530);
   U2862 : aoi12 port map( b => n1973, c => n1971, a => n1974, outb => n1970);
   U2863 : nand3 port map( a => n1975, b => n1976, c => n1977, outb => 
                           display_out_n529);
   U2864 : nand2 port map( a => n1978, b => n1972, outb => n1977);
   U2865 : nand2 port map( a => display_out_clk_timer_4_port, b => n231, outb 
                           => n1976);
   U2866 : oai12 port map( b => n230, c => n226, a => n1972, outb => n231);
   U2867 : nand3 port map( a => n230, b => n222, c => n229, outb => n1975);
   U2868 : inv port map( inb => display_out_clk_timer_4_port, outb => n229);
   U2869 : inv port map( inb => n1979, outb => n230);
   U2870 : oai22 port map( a => n1980, b => n235, c => n1981, d => n1972, outb 
                           => display_out_n528);
   U2871 : aoi12 port map( b => n1973, c => n1982, a => n1974, outb => n1980);
   U2872 : oai12 port map( b => n1983, c => n1981, a => n1979, outb => n1982);
   U2873 : oai12 port map( b => n235, c => n1984, a => n1985, outb => 
                           display_out_n527);
   U2874 : aoi22 port map( a => display_out_clk_timer_2_port, b => n1986, c => 
                           n1983, d => n222, outb => n1985);
   U2875 : inv port map( inb => n226, outb => n222);
   U2876 : oai12 port map( b => n1987, c => n226, a => n1972, outb => n1986);
   U2877 : nor2 port map( a => n1988, b => n1989, outb => n226);
   U2878 : inv port map( inb => n1972, outb => n235);
   U2879 : nand4 port map( a => n1990, b => n1991, c => n1992, d => n1993, outb
                           => n1972);
   U2880 : nand2 port map( a => n1994, b => n1942, outb => n1992);
   U2881 : inv port map( inb => n1995, outb => n1942);
   U2882 : inv port map( inb => n1988, outb => n1991);
   U2883 : nand2 port map( a => n1996, b => n1997, outb => n1988);
   U2884 : nand2 port map( a => n1998, b => n1999, outb => display_out_n526);
   U2885 : aoi22 port map( a => n248, b => n2000, c => n256, d => 
                           display_out_disp_timer_0_port, outb => n1998);
   U2886 : nand3 port map( a => n2001, b => n2002, c => n2003, outb => 
                           display_out_n525);
   U2887 : nand2 port map( a => n303, b => n248, outb => n2003);
   U2888 : oai12 port map( b => n2004, c => n2005, a => 
                           display_out_disp_timer_15_port, outb => n2001);
   U2889 : nor2 port map( a => n244, b => n2006, outb => n2004);
   U2890 : nand4 port map( a => n2007, b => n2002, c => n2008, d => n2009, outb
                           => display_out_n524);
   U2891 : nand2 port map( a => display_out_disp_timer_14_port, b => n2005, 
                           outb => n2009);
   U2892 : oai12 port map( b => n244, c => n2010, a => n265, outb => n2005);
   U2893 : nand3 port map( a => n2010, b => n248, c => n2006, outb => n2008);
   U2894 : nand3 port map( a => n2011, b => n2007, c => n2012, outb => 
                           display_out_n523);
   U2895 : aoi22 port map( a => display_out_disp_timer_13_port, b => n2013, c 
                           => n2010, d => n248, outb => n2012);
   U2896 : inv port map( inb => n2014, outb => n2010);
   U2897 : inv port map( inb => n2015, outb => n2013);
   U2898 : aoi12 port map( b => n248, c => display_out_disp_timer_12_port, a =>
                           n2016, outb => n2015);
   U2899 : nand4 port map( a => n2011, b => n2017, c => n2018, d => n2019, outb
                           => display_out_n522);
   U2900 : nand2 port map( a => display_out_disp_timer_12_port, b => n2016, 
                           outb => n2019);
   U2901 : oai12 port map( b => n244, c => n2020, a => n265, outb => n2016);
   U2902 : nand3 port map( a => n2020, b => n248, c => n2021, outb => n2018);
   U2903 : nand4 port map( a => n2017, b => n2002, c => n2022, d => n2023, outb
                           => display_out_n521);
   U2904 : aoi22 port map( a => display_out_disp_timer_11_port, b => n2024, c 
                           => n2020, d => n248, outb => n2023);
   U2905 : nand2 port map( a => n265, b => n2025, outb => n2024);
   U2906 : oai12 port map( b => display_out_disp_timer_10_port, c => n2026, a 
                           => n248, outb => n2025);
   U2907 : nand3 port map( a => n2027, b => display_out_bcd_time_2_port, c => 
                           n2028, outb => n2017);
   U2908 : inv port map( inb => n2029, outb => n2027);
   U2909 : nand4 port map( a => n2030, b => n2002, c => n2031, d => n2032, outb
                           => display_out_n520);
   U2910 : oai12 port map( b => n2033, c => n256, a => 
                           display_out_disp_timer_10_port, outb => n2032);
   U2911 : nor2 port map( a => n244, b => n2034, outb => n2033);
   U2912 : inv port map( inb => n2035, outb => n2031);
   U2913 : nor3 port map( a => n2026, b => n244, c => 
                           display_out_disp_timer_10_port, outb => n2035);
   U2914 : nand2 port map( a => n1959, b => n2028, outb => n2002);
   U2915 : nor3 port map( a => display_out_bcd_time_1_port, b => 
                           display_out_bcd_time_2_port, c => 
                           display_out_bcd_time_0_port, outb => n1959);
   U2916 : inv port map( inb => n2036, outb => n2030);
   U2917 : nor2 port map( a => n2037, b => n2038, outb => n2036);
   U2918 : nand3 port map( a => n2039, b => n2007, c => n2040, outb => 
                           display_out_n519);
   U2919 : aoi22 port map( a => n2028, b => n2041, c => n2034, d => n248, outb 
                           => n2040);
   U2920 : inv port map( inb => n2026, outb => n2034);
   U2921 : nand2 port map( a => n2042, b => n2028, outb => n2007);
   U2922 : oai12 port map( b => n2043, c => n2044, a => 
                           display_out_disp_timer_9_port, outb => n2039);
   U2923 : nor2 port map( a => n244, b => n2045, outb => n2043);
   U2924 : nand4 port map( a => n2046, b => n2011, c => n2047, d => n2048, outb
                           => display_out_n518);
   U2925 : nand2 port map( a => display_out_disp_timer_8_port, b => n2044, outb
                           => n2048);
   U2926 : oai12 port map( b => n244, c => n2049, a => n265, outb => n2044);
   U2927 : nand3 port map( a => n2049, b => n248, c => n2045, outb => n2047);
   U2928 : nand2 port map( a => n2050, b => n2028, outb => n2011);
   U2929 : nand3 port map( a => n2051, b => n2022, c => n2052, outb => 
                           display_out_n517);
   U2930 : aoi22 port map( a => n2049, b => n248, c => n2053, d => n265, outb 
                           => n2052);
   U2931 : oai12 port map( b => n256, c => n2054, a => 
                           display_out_disp_timer_7_port, outb => n2051);
   U2932 : oai12 port map( b => n2038, c => n2037, a => n2055, outb => 
                           display_out_n516);
   U2933 : inv port map( inb => n2056, outb => n2055);
   U2934 : oai22 port map( a => n2057, b => n2058, c => n2054, d => n244, outb 
                           => n2056);
   U2935 : aoi12 port map( b => n248, c => display_out_disp_timer_5_port, a => 
                           n2059, outb => n2058);
   U2936 : nor3 port map( a => n2060, b => n2042, c => n2061, outb => n2038);
   U2937 : nand3 port map( a => n2062, b => n2063, c => n2064, outb => 
                           display_out_n515);
   U2938 : nand2 port map( a => n2028, b => n2041, outb => n2064);
   U2939 : inv port map( inb => n2065, outb => n2041);
   U2940 : nor3 port map( a => n2050, b => n2066, c => n2061, outb => n2065);
   U2941 : nor3 port map( a => n2067, b => display_out_bcd_time_0_port, c => 
                           n1956, outb => n2050);
   U2942 : nand2 port map( a => display_out_disp_timer_5_port, b => n2059, outb
                           => n2063);
   U2943 : oai12 port map( b => n244, c => n2068, a => n265, outb => n2059);
   U2944 : nand3 port map( a => n2068, b => n248, c => n2069, outb => n2062);
   U2945 : nand2 port map( a => n2070, b => n2046, outb => display_out_n514);
   U2946 : aoi22 port map( a => n2028, b => n2066, c => n265, d => n2053, outb 
                           => n2046);
   U2947 : oai12 port map( b => n2071, c => n2029, a => n2072, outb => n2053);
   U2948 : aoi22 port map( a => display_out_disp_timer_4_port, b => n2073, c =>
                           n2068, d => n248, outb => n2070);
   U2949 : nand3 port map( a => n265, b => n2074, c => n2075, outb => n2073);
   U2950 : nand4 port map( a => n1999, b => n2022, c => n2076, d => n2077, outb
                           => display_out_n513);
   U2951 : oai12 port map( b => n256, c => n2078, a => 
                           display_out_disp_timer_3_port, outb => n2077);
   U2952 : inv port map( inb => n265, outb => n256);
   U2953 : nand3 port map( a => n2075, b => n248, c => n2074, outb => n2076);
   U2954 : nand2 port map( a => n2060, b => n2028, outb => n2022);
   U2955 : inv port map( inb => n2037, outb => n2028);
   U2956 : nor3 port map( a => display_out_bcd_time_0_port, b => 
                           display_out_bcd_time_1_port, c => n1956, outb => 
                           n2060);
   U2957 : nor2 port map( a => n1974, b => n2079, outb => n1999);
   U2958 : nor3 port map( a => n2029, b => display_out_bcd_time_2_port, c => 
                           n2037, outb => n2079);
   U2959 : nand2 port map( a => display_out_bcd_time_0_port, b => n2067, outb 
                           => n2029);
   U2960 : oai12 port map( b => n2037, c => n2080, a => n2081, outb => 
                           display_out_n512);
   U2961 : aoi22 port map( a => display_out_disp_timer_2_port, b => n2082, c =>
                           n2075, d => n248, outb => n2081);
   U2962 : oai12 port map( b => n244, c => n2083, a => n265, outb => n2082);
   U2963 : inv port map( inb => n2061, outb => n2080);
   U2964 : nor3 port map( a => n2084, b => display_out_bcd_time_2_port, c => 
                           n2067, outb => n2061);
   U2965 : oai12 port map( b => n2037, c => n2085, a => n2086, outb => 
                           display_out_n511);
   U2966 : aoi22 port map( a => display_out_disp_timer_1_port, b => n2087, c =>
                           n2083, d => n248, outb => n2086);
   U2967 : inv port map( inb => n244, outb => n248);
   U2968 : oai12 port map( b => n244, c => n2000, a => n265, outb => n2087);
   U2969 : inv port map( inb => display_out_disp_timer_0_port, outb => n2000);
   U2970 : nor2 port map( a => n1973, b => n1965, outb => n244);
   U2971 : nand3 port map( a => n1949, b => n1996, c => n1993, outb => n1973);
   U2972 : inv port map( inb => n2066, outb => n2085);
   U2973 : nor3 port map( a => display_out_bcd_time_0_port, b => 
                           display_out_bcd_time_2_port, c => n2067, outb => 
                           n2066);
   U2974 : nand2 port map( a => n1947, b => n265, outb => n2037);
   U2975 : nand4 port map( a => n1966, b => n2088, c => n1993, d => n1996, outb
                           => n265);
   U2976 : aoi12 port map( b => n1978, c => n2089, a => n1965, outb => n1966);
   U2977 : nor2 port map( a => n2090, b => n1984, outb => n1965);
   U2978 : oai22 port map( a => n1955, b => n2084, c => n2091, d => n1958, outb
                           => display_out_n510);
   U2979 : oai22 port map( a => n1955, b => n2067, c => n1951, d => n1958, outb
                           => display_out_n509);
   U2980 : xor2 port map( a => n1947, b => n2092, outb => n1951);
   U2981 : oai12 port map( b => n2093, c => n2094, a => n2095, outb => 
                           display_out_n508);
   U2982 : nand2 port map( a => hub_blank_o_port, b => n2094, outb => n2095);
   U2983 : nor2 port map( a => n2096, b => n1994, outb => n2094);
   U2984 : inv port map( inb => n1967, outb => n1994);
   U2985 : nor2 port map( a => n1978, b => n1974, outb => n2093);
   U2986 : nand2 port map( a => n2072, b => n2097, outb => display_out_n507);
   U2987 : nand2 port map( a => hub_mux_o_2_port, b => n2098, outb => n2097);
   U2988 : inv port map( inb => n2099, outb => display_out_n506);
   U2989 : aoi22 port map( a => n2098, b => display_out_h_row_0_port, c => 
                           n2100, d => n2101, outb => n2099);
   U2990 : oai12 port map( b => n2102, c => n2103, a => n2104, outb => 
                           display_out_n505);
   U2991 : nand3 port map( a => n2101, b => display_out_h_row_0_port, c => 
                           n2103, outb => n2104);
   U2992 : inv port map( inb => display_out_h_row_1_port, outb => n2103);
   U2993 : aoi12 port map( b => n1978, c => n2100, a => n2098, outb => n2102);
   U2994 : inv port map( inb => display_out_h_row_0_port, outb => n2100);
   U2995 : nand3 port map( a => n2105, b => n2072, c => n2106, outb => 
                           display_out_n504);
   U2996 : nand2 port map( a => hub_mux_o_0_port, b => n2098, outb => n2106);
   U2997 : nand2 port map( a => n2101, b => display_out_h_row_0_port, outb => 
                           n2105);
   U2998 : nand3 port map( a => n2107, b => n2072, c => n2108, outb => 
                           display_out_n503);
   U2999 : nand2 port map( a => hub_mux_o_1_port, b => n2098, outb => n2108);
   U3000 : nand2 port map( a => display_out_h_row_1_port, b => n2101, outb => 
                           n2107);
   U3001 : nor2 port map( a => n1984, b => n2098, outb => n2101);
   U3002 : inv port map( inb => n2096, outb => n2098);
   U3003 : nand2 port map( a => n2072, b => n2109, outb => n2096);
   U3004 : nand3 port map( a => n1947, b => n2089, c => n2042, outb => n2109);
   U3005 : nor3 port map( a => n2067, b => n2084, c => n1956, outb => n2042);
   U3006 : inv port map( inb => display_out_bcd_time_0_port, outb => n2084);
   U3007 : inv port map( inb => n245, outb => n2089);
   U3008 : nand2 port map( a => n1962, b => n2110, outb => display_out_n502);
   U3009 : nand3 port map( a => n1968, b => n1984, c => hub_clk_o_port, outb =>
                           n2110);
   U3010 : nor3 port map( a => n1974, b => n2111, c => n1969, outb => n1968);
   U3011 : aoi12 port map( b => n1941, c => n2111, a => n1989, outb => n1962);
   U3012 : nor2 port map( a => n1993, b => n223, outb => n1989);
   U3013 : inv port map( inb => n1996, outb => n2111);
   U3014 : oai22 port map( a => n2112, b => n2113, c => n59, d => n2114, outb 
                           => display_out_n501);
   U3015 : inv port map( inb => n2113, outb => n2114);
   U3016 : inv port map( inb => hub_reg_f, outb => n59);
   U3017 : nor2 port map( a => n2115, b => n1937, outb => n2113);
   U3018 : nor2 port map( a => n1996, b => n1941, outb => n1937);
   U3019 : inv port map( inb => n2116, outb => n1941);
   U3020 : inv port map( inb => n2117, outb => n2115);
   U3021 : nor2 port map( a => n1939, b => n1943, outb => n2112);
   U3022 : oai22 port map( a => n2091, b => n1952, c => n2118, d => n1954, outb
                           => display_out_n500);
   U3023 : oai22 port map( a => n1961, b => n1952, c => n2119, d => n1954, outb
                           => display_out_n499);
   U3024 : nand2 port map( a => n1969, b => n1954, outb => n1952);
   U3025 : nand2 port map( a => n2117, b => n2120, outb => n1954);
   U3026 : nor2 port map( a => n2121, b => n1974, outb => n2117);
   U3027 : aoi22 port map( a => n2122, b => n2123, c => n2071, d => n2124, outb
                           => n1961);
   U3028 : inv port map( inb => n2125, outb => n2124);
   U3029 : nand3 port map( a => n1947, b => n2125, c => n2092, outb => n2123);
   U3030 : oai12 port map( b => n2126, c => n2091, a => n2125, outb => n2092);
   U3031 : nand2 port map( a => n2126, b => n2091, outb => n2125);
   U3032 : inv port map( inb => n2127, outb => n2091);
   U3033 : aoi12 port map( b => n1947, c => display_out_bcd_time_0_port, a => 
                           n2128, outb => n2127);
   U3034 : oai12 port map( b => n2071, c => n2067, a => n2129, outb => n2126);
   U3035 : inv port map( inb => display_out_bcd_time_1_port, outb => n2067);
   U3036 : inv port map( inb => n2071, outb => n1947);
   U3037 : oai22 port map( a => n1956, b => n2071, c => n2120, d => n2119, outb
                           => n2122);
   U3038 : inv port map( inb => display_out_h_col_2_port, outb => n2119);
   U3039 : inv port map( inb => display_out_bcd_time_2_port, outb => n1956);
   U3040 : nand3 port map( a => n1958, b => n1997, c => n2130, outb => 
                           display_out_n498);
   U3041 : nand3 port map( a => n1990, b => n1967, c => hub_latch_o_port, outb 
                           => n2130);
   U3042 : nand2 port map( a => n1943, b => n223, outb => n1967);
   U3043 : inv port map( inb => n1955, outb => n1990);
   U3044 : nand2 port map( a => n1943, b => n2116, outb => n1997);
   U3045 : nand2 port map( a => n1978, b => n1955, outb => n1958);
   U3046 : oai12 port map( b => n245, c => n2071, a => n2072, outb => n1955);
   U3047 : nand2 port map( a => n1978, b => n2090, outb => n2071);
   U3048 : nand2 port map( a => n2131, b => n247, outb => n2090);
   U3049 : nand3 port map( a => n2132, b => n2133, c => n2134, outb => n2131);
   U3050 : nor3 port map( a => n2135, b => n2136, c => n2137, outb => n2134);
   U3051 : nand4 port map( a => n2138, b => n2074, c => n2139, d => n2069, outb
                           => n2137);
   U3052 : inv port map( inb => display_out_disp_timer_4_port, outb => n2139);
   U3053 : inv port map( inb => display_out_disp_timer_3_port, outb => n2074);
   U3054 : nand4 port map( a => n2057, b => n2140, c => n2045, d => n2141, outb
                           => n2136);
   U3055 : inv port map( inb => display_out_disp_timer_7_port, outb => n2140);
   U3056 : nand4 port map( a => n262, b => n258, c => n2142, d => n2143, outb 
                           => n2135);
   U3057 : nor3 port map( a => display_out_disp_timer_24_port, b => 
                           display_out_disp_timer_26_port, c => 
                           display_out_disp_timer_25_port, outb => n2143);
   U3058 : nor2 port map( a => display_out_disp_timer_2_port, b => 
                           display_out_disp_timer_29_port, outb => n2142);
   U3059 : nor2 port map( a => n2144, b => n2145, outb => n2133);
   U3060 : nand4 port map( a => n301, b => n298, c => n292, d => n2146, outb =>
                           n2145);
   U3061 : nand4 port map( a => n285, b => n2147, c => n280, d => n277, outb =>
                           n2144);
   U3062 : inv port map( inb => display_out_disp_timer_21_port, outb => n2147);
   U3063 : inv port map( inb => display_out_disp_timer_20_port, outb => n285);
   U3064 : nor3 port map( a => n2148, b => n2149, c => n2150, outb => n2132);
   U3065 : inv port map( inb => n2151, outb => n2150);
   U3066 : nor2 port map( a => display_out_disp_timer_10_port, b => 
                           display_out_disp_timer_11_port, outb => n2151);
   U3067 : nand4 port map( a => n2021, b => n2152, c => n2006, d => n2153, outb
                           => n2148);
   U3068 : inv port map( inb => display_out_disp_timer_15_port, outb => n2153);
   U3069 : inv port map( inb => display_out_disp_timer_14_port, outb => n2006);
   U3070 : nand4 port map( a => n259, b => n253, c => n2138, d => n247, outb =>
                           n245);
   U3071 : inv port map( inb => display_out_disp_timer_31_port, outb => n247);
   U3072 : inv port map( inb => display_out_disp_timer_30_port, outb => n2138);
   U3073 : inv port map( inb => display_out_disp_timer_29_port, outb => n253);
   U3074 : inv port map( inb => n255, outb => n259);
   U3075 : nand3 port map( a => n262, b => n258, c => n264, outb => n255);
   U3076 : nor3 port map( a => display_out_disp_timer_25_port, b => 
                           display_out_disp_timer_26_port, c => n2154, outb => 
                           n264);
   U3077 : inv port map( inb => n271, outb => n2154);
   U3078 : nor2 port map( a => n275, b => display_out_disp_timer_24_port, outb 
                           => n271);
   U3079 : nand3 port map( a => n280, b => n277, c => n282, outb => n275);
   U3080 : nor3 port map( a => display_out_disp_timer_20_port, b => 
                           display_out_disp_timer_21_port, c => n289, outb => 
                           n282);
   U3081 : nand3 port map( a => n292, b => n2146, c => n295, outb => n289);
   U3082 : inv port map( inb => n296, outb => n295);
   U3083 : nand3 port map( a => n301, b => n298, c => n303, outb => n296);
   U3084 : nor3 port map( a => display_out_disp_timer_14_port, b => 
                           display_out_disp_timer_15_port, c => n2014, outb => 
                           n303);
   U3085 : nand3 port map( a => n2021, b => n2152, c => n2020, outb => n2014);
   U3086 : nor3 port map( a => display_out_disp_timer_10_port, b => 
                           display_out_disp_timer_11_port, c => n2026, outb => 
                           n2020);
   U3087 : nand3 port map( a => n2045, b => n2141, c => n2049, outb => n2026);
   U3088 : nor2 port map( a => n2054, b => display_out_disp_timer_7_port, outb 
                           => n2049);
   U3089 : nand3 port map( a => n2069, b => n2057, c => n2068, outb => n2054);
   U3090 : nor3 port map( a => display_out_disp_timer_3_port, b => 
                           display_out_disp_timer_4_port, c => n2078, outb => 
                           n2068);
   U3091 : inv port map( inb => n2075, outb => n2078);
   U3092 : nor2 port map( a => n2149, b => display_out_disp_timer_2_port, outb 
                           => n2075);
   U3093 : inv port map( inb => n2083, outb => n2149);
   U3094 : nor2 port map( a => display_out_disp_timer_1_port, b => 
                           display_out_disp_timer_0_port, outb => n2083);
   U3095 : inv port map( inb => display_out_disp_timer_6_port, outb => n2057);
   U3096 : inv port map( inb => display_out_disp_timer_5_port, outb => n2069);
   U3097 : inv port map( inb => display_out_disp_timer_9_port, outb => n2141);
   U3098 : inv port map( inb => display_out_disp_timer_8_port, outb => n2045);
   U3099 : inv port map( inb => display_out_disp_timer_13_port, outb => n2152);
   U3100 : inv port map( inb => display_out_disp_timer_12_port, outb => n2021);
   U3101 : inv port map( inb => display_out_disp_timer_17_port, outb => n298);
   U3102 : inv port map( inb => display_out_disp_timer_16_port, outb => n301);
   U3103 : inv port map( inb => display_out_disp_timer_19_port, outb => n2146);
   U3104 : inv port map( inb => display_out_disp_timer_18_port, outb => n292);
   U3105 : inv port map( inb => display_out_disp_timer_23_port, outb => n277);
   U3106 : inv port map( inb => display_out_disp_timer_22_port, outb => n280);
   U3107 : inv port map( inb => display_out_disp_timer_28_port, outb => n258);
   U3108 : inv port map( inb => display_out_disp_timer_27_port, outb => n262);
   U3109 : inv port map( inb => n1984, outb => n1978);
   U3110 : nand3 port map( a => display_out_hub_out_sm_0_port, b => n1945, c =>
                           display_out_hub_out_sm_1_port, outb => n1984);
   U3111 : oai12 port map( b => n2155, c => n2156, a => n2157, outb => 
                           display_out_n497);
   U3112 : aoi22 port map( a => display_out_hub_piso_r0_2_port, b => n2158, c 
                           => n2159, d => mem_sipo_r0_1_port, outb => n2157);
   U3113 : inv port map( inb => display_out_hub_piso_r0_1_port, outb => n2156);
   U3114 : oai12 port map( b => n2160, c => n2155, a => n2161, outb => 
                           display_out_n496);
   U3115 : aoi22 port map( a => display_out_hub_piso_r0_3_port, b => n2158, c 
                           => n2159, d => mem_sipo_r0_2_port, outb => n2161);
   U3116 : inv port map( inb => display_out_hub_piso_r0_2_port, outb => n2160);
   U3117 : oai12 port map( b => n2155, c => n2162, a => n2163, outb => 
                           display_out_n495);
   U3118 : aoi22 port map( a => display_out_hub_piso_r0_4_port, b => n2158, c 
                           => n2159, d => mem_sipo_r0_3_port, outb => n2163);
   U3119 : inv port map( inb => display_out_hub_piso_r0_3_port, outb => n2162);
   U3120 : oai12 port map( b => n2155, c => n2164, a => n2165, outb => 
                           display_out_n494);
   U3121 : aoi22 port map( a => display_out_hub_piso_r0_5_port, b => n2158, c 
                           => n2159, d => mem_sipo_r0_4_port, outb => n2165);
   U3122 : inv port map( inb => display_out_hub_piso_r0_4_port, outb => n2164);
   U3123 : oai12 port map( b => n2155, c => n2166, a => n2167, outb => 
                           display_out_n493);
   U3124 : aoi22 port map( a => display_out_hub_piso_r0_6_port, b => n2158, c 
                           => n2159, d => mem_sipo_r0_5_port, outb => n2167);
   U3125 : inv port map( inb => display_out_hub_piso_r0_5_port, outb => n2166);
   U3126 : oai12 port map( b => n2155, c => n2168, a => n2169, outb => 
                           display_out_n492);
   U3127 : aoi22 port map( a => n2158, b => display_out_hub_piso_r0_7_port, c 
                           => n2159, d => mem_sipo_r0_6_port, outb => n2169);
   U3128 : inv port map( inb => display_out_hub_piso_r0_6_port, outb => n2168);
   U3129 : oai12 port map( b => n2155, c => n2170, a => n2171, outb => 
                           display_out_n491);
   U3130 : aoi22 port map( a => display_out_hub_piso_r0_1_port, b => n2158, c 
                           => n2159, d => mem_sipo_r0_0_port, outb => n2171);
   U3131 : oai12 port map( b => n2155, c => n2172, a => n2173, outb => 
                           display_out_n490);
   U3132 : aoi22 port map( a => display_out_hub_piso_g0_2_port, b => n2158, c 
                           => n2159, d => mem_sipo_g0_1_port, outb => n2173);
   U3133 : inv port map( inb => display_out_hub_piso_g0_1_port, outb => n2172);
   U3134 : oai12 port map( b => n2155, c => n2174, a => n2175, outb => 
                           display_out_n489);
   U3135 : aoi22 port map( a => display_out_hub_piso_g0_3_port, b => n2158, c 
                           => n2159, d => mem_sipo_g0_2_port, outb => n2175);
   U3136 : inv port map( inb => display_out_hub_piso_g0_2_port, outb => n2174);
   U3137 : oai12 port map( b => n2155, c => n2176, a => n2177, outb => 
                           display_out_n488);
   U3138 : aoi22 port map( a => display_out_hub_piso_g0_4_port, b => n2158, c 
                           => n2159, d => mem_sipo_g0_3_port, outb => n2177);
   U3139 : inv port map( inb => display_out_hub_piso_g0_3_port, outb => n2176);
   U3140 : oai12 port map( b => n2155, c => n2178, a => n2179, outb => 
                           display_out_n487);
   U3141 : aoi22 port map( a => display_out_hub_piso_g0_5_port, b => n2158, c 
                           => n2159, d => mem_sipo_g0_4_port, outb => n2179);
   U3142 : inv port map( inb => display_out_hub_piso_g0_4_port, outb => n2178);
   U3143 : oai12 port map( b => n2155, c => n2180, a => n2181, outb => 
                           display_out_n486);
   U3144 : aoi22 port map( a => display_out_hub_piso_g0_6_port, b => n2158, c 
                           => n2159, d => mem_sipo_g0_5_port, outb => n2181);
   U3145 : inv port map( inb => display_out_hub_piso_g0_5_port, outb => n2180);
   U3146 : oai12 port map( b => n2155, c => n2182, a => n2183, outb => 
                           display_out_n485);
   U3147 : aoi22 port map( a => n2158, b => display_out_hub_piso_g0_7_port, c 
                           => n2159, d => mem_sipo_g0_6_port, outb => n2183);
   U3148 : inv port map( inb => display_out_hub_piso_g0_6_port, outb => n2182);
   U3149 : oai12 port map( b => n2155, c => n2184, a => n2185, outb => 
                           display_out_n484);
   U3150 : aoi22 port map( a => display_out_hub_piso_g0_1_port, b => n2158, c 
                           => n2159, d => mem_sipo_g0_0_port, outb => n2185);
   U3151 : oai12 port map( b => n2155, c => n2186, a => n2187, outb => 
                           display_out_n483);
   U3152 : aoi22 port map( a => display_out_hub_piso_b0_2_port, b => n2158, c 
                           => n2159, d => mem_sipo_b0_1_port, outb => n2187);
   U3153 : inv port map( inb => display_out_hub_piso_b0_1_port, outb => n2186);
   U3154 : oai12 port map( b => n2155, c => n2188, a => n2189, outb => 
                           display_out_n482);
   U3155 : aoi22 port map( a => display_out_hub_piso_b0_3_port, b => n2158, c 
                           => n2159, d => mem_sipo_b0_2_port, outb => n2189);
   U3156 : inv port map( inb => display_out_hub_piso_b0_2_port, outb => n2188);
   U3157 : oai12 port map( b => n2155, c => n2190, a => n2191, outb => 
                           display_out_n481);
   U3158 : aoi22 port map( a => display_out_hub_piso_b0_4_port, b => n2158, c 
                           => n2159, d => mem_sipo_b0_3_port, outb => n2191);
   U3159 : inv port map( inb => display_out_hub_piso_b0_3_port, outb => n2190);
   U3160 : oai12 port map( b => n2155, c => n2192, a => n2193, outb => 
                           display_out_n480);
   U3161 : aoi22 port map( a => display_out_hub_piso_b0_5_port, b => n2158, c 
                           => n2159, d => mem_sipo_b0_4_port, outb => n2193);
   U3162 : inv port map( inb => display_out_hub_piso_b0_4_port, outb => n2192);
   U3163 : oai12 port map( b => n2155, c => n2194, a => n2195, outb => 
                           display_out_n479);
   U3164 : aoi22 port map( a => display_out_hub_piso_b0_6_port, b => n2158, c 
                           => n2159, d => mem_sipo_b0_5_port, outb => n2195);
   U3165 : inv port map( inb => display_out_hub_piso_b0_5_port, outb => n2194);
   U3166 : oai12 port map( b => n2155, c => n2196, a => n2197, outb => 
                           display_out_n478);
   U3167 : aoi22 port map( a => n2158, b => display_out_hub_piso_b0_7_port, c 
                           => n2159, d => mem_sipo_b0_6_port, outb => n2197);
   U3168 : inv port map( inb => display_out_hub_piso_b0_6_port, outb => n2196);
   U3169 : oai12 port map( b => n2155, c => n2198, a => n2199, outb => 
                           display_out_n477);
   U3170 : aoi22 port map( a => display_out_hub_piso_b0_1_port, b => n2158, c 
                           => n2159, d => mem_sipo_b0_0_port, outb => n2199);
   U3171 : nor2 port map( a => n2088, b => n2200, outb => n2159);
   U3172 : nor2 port map( a => n1943, b => n1974, outb => n2088);
   U3173 : inv port map( inb => n2072, outb => n1974);
   U3174 : inv port map( inb => n1949, outb => n1943);
   U3175 : nor2 port map( a => n1993, b => n2200, outb => n2158);
   U3176 : inv port map( inb => n2155, outb => n2200);
   U3177 : nand2 port map( a => n217, b => n2120, outb => n2155);
   U3178 : nand2 port map( a => n1938, b => n2116, outb => n2120);
   U3179 : nor2 port map( a => n2121, b => n1939, outb => n217);
   U3180 : nor2 port map( a => n2072, b => n1995, outb => n1939);
   U3181 : nand3 port map( a => n2201, b => n1945, c => n2202, outb => n2072);
   U3182 : nor3 port map( a => n2116, b => n1995, c => n1949, outb => n2121);
   U3183 : nand3 port map( a => n2202, b => n2201, c => 
                           display_out_hub_out_sm_2_port, outb => n1949);
   U3184 : nand2 port map( a => mem_hub_f, b => reg_hub_f, outb => n1995);
   U3185 : nand4 port map( a => n2203, b => n2204, c => n2205, d => n1981, outb
                           => n2116);
   U3186 : nand3 port map( a => n2206, b => n1996, c => n2207, outb => n2205);
   U3187 : nand2 port map( a => n2208, b => n2209, outb => n2207);
   U3188 : nand2 port map( a => display_out_h_col_2_port, b => n1938, outb => 
                           n2206);
   U3189 : inv port map( inb => n2210, outb => n2204);
   U3190 : nor2 port map( a => n2209, b => n2208, outb => n2210);
   U3191 : nor2 port map( a => n1938, b => display_out_clk_timer_2_port, outb 
                           => n2208);
   U3192 : oai22 port map( a => n2211, b => n2129, c => n2211, d => n2212, outb
                           => n2209);
   U3193 : nand2 port map( a => n2213, b => n234, outb => n2212);
   U3194 : inv port map( inb => display_out_clk_timer_1_port, outb => n234);
   U3195 : nand2 port map( a => display_out_h_col_1_port, b => n1938, outb => 
                           n2129);
   U3196 : inv port map( inb => n2213, outb => n1938);
   U3197 : aoi12 port map( b => n1971, c => n2213, a => n2128, outb => n2211);
   U3198 : nor2 port map( a => n2118, b => n2213, outb => n2128);
   U3199 : inv port map( inb => display_out_h_col_0_port, outb => n2118);
   U3200 : nand2 port map( a => n223, b => n1969, outb => n2213);
   U3201 : inv port map( inb => n1993, outb => n1969);
   U3202 : nand3 port map( a => n2202, b => n1945, c => 
                           display_out_hub_out_sm_1_port, outb => n1993);
   U3203 : inv port map( inb => display_out_hub_out_sm_0_port, outb => n2202);
   U3204 : nor2 port map( a => n1979, b => n2214, outb => n223);
   U3205 : inv port map( inb => n2203, outb => n2214);
   U3206 : nand2 port map( a => n1983, b => n1981, outb => n1979);
   U3207 : inv port map( inb => display_out_clk_timer_3_port, outb => n1981);
   U3208 : nor2 port map( a => n232, b => display_out_clk_timer_2_port, outb =>
                           n1983);
   U3209 : inv port map( inb => n1987, outb => n232);
   U3210 : nor2 port map( a => display_out_clk_timer_0_port, b => 
                           display_out_clk_timer_1_port, outb => n1987);
   U3211 : inv port map( inb => display_out_clk_timer_0_port, outb => n1971);
   U3212 : nor3 port map( a => display_out_clk_timer_5_port, b => 
                           display_out_clk_timer_6_port, c => 
                           display_out_clk_timer_4_port, outb => n2203);
   U3213 : oai12 port map( b => n1996, c => n2170, a => n2215, outb => 
                           display_out_n476);
   U3214 : nand2 port map( a => hub_r0_o_port, b => n1996, outb => n2215);
   U3215 : inv port map( inb => display_out_hub_piso_r0_0_port, outb => n2170);
   U3216 : oai12 port map( b => n1996, c => n2184, a => n2216, outb => 
                           display_out_n475);
   U3217 : nand2 port map( a => hub_g0_o_port, b => n1996, outb => n2216);
   U3218 : inv port map( inb => display_out_hub_piso_g0_0_port, outb => n2184);
   U3219 : oai12 port map( b => n1996, c => n2198, a => n2217, outb => 
                           display_out_n474);
   U3220 : nand2 port map( a => hub_b0_o_port, b => n1996, outb => n2217);
   U3221 : inv port map( inb => display_out_hub_piso_b0_0_port, outb => n2198);
   U3222 : nand3 port map( a => n2201, b => n1945, c => 
                           display_out_hub_out_sm_0_port, outb => n1996);
   U3223 : inv port map( inb => display_out_hub_out_sm_2_port, outb => n1945);
   U3224 : inv port map( inb => display_out_hub_out_sm_1_port, outb => n2201);

end SYN_rtl;
