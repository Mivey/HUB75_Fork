library IEEE;
use IEEE.std_logic_1164.all;

entity inv is
port(a: in STD_logic;
     b: out STD_Logic);
end inv;
architecture structure of inv is
begin
b <= not (a);
end structure;

library IEEE;
use IEEE.std_logic_1164.all;

entity nand2 is
port(a, b: in STD_logic;
	c: out STD_Logic);
end nand2;
architecture structure of nand2 is
begin
c <= not(a and b);
end structure;

library IEEE;
use IEEE.std_logic_1164.all;

entity nand3 is
port(a, b, c: in STD_logic;
           d: out STD_Logic);
end nand3 ;
architecture structure of nand3 is
begin
d <= not(a and b and c);
end structure;

library IEEE;
use IEEE.std_logic_1164.all;

entity nand4 is
port(a, b, c, d: in STD_logic;
	      e: out STD_Logic);
end nand4 ;
architecture structure of nand4 is
begin
e <= not(a and b and c and d);
end structure;

library IEEE;
use IEEE.std_logic_1164.all;

entity nor2 is
port(a, b: in STD_logic;
	c: out STD_Logic);
end nor2 ;
architecture structure of nor2 is
begin
c <= not(a or b);
end structure;

library IEEE;
use IEEE.std_logic_1164.all;

entity nor3 is
port(a, b, c: in STD_logic;
	   d: out STD_Logic);
end nor3 ;
architecture structure of nor3 is
begin
d <= not(a or b or c);
end structure;

library IEEE;
use IEEE.std_logic_1164.all;

entity xor2 is
port(a, b: in STD_logic;
        c: out STD_Logic);
end xor2 ;
architecture structure of xor2 is
begin
c <= (a xor b);
end structure;

library IEEE;
use IEEE.std_logic_1164.all;

entity aoi12 is
port(a, b, c: in STD_logic;
	   d: out STD_Logic);
end aoi12 ;
architecture structure of aoi12 is
begin
d <= not(a or (b and c));
end structure;

library IEEE;
use IEEE.std_logic_1164.all;

entity aoi22 is
port(a, b, c, d: in STD_logic;
              e: out STD_Logic);
end aoi22 ;
architecture structure of aoi22 is
begin
e <= not((a and b) or (c and d));
end structure;


library IEEE;
use IEEE.std_logic_1164.all;

entity oai12 is
port(a, b, c: in STD_logic;
	   d: out STD_Logic);
end oai12;
architecture structure of oai12 is
begin
d <= not(a and (b or c));
end structure;

library IEEE;
use IEEE.std_logic_1164.all;

entity oai22 is
port(a, b, c, d: in STD_logic;
              e: out STD_Logic);
end oai22; 
architecture structure of oai22 is
begin
e <= not((a or b) and (c or d));
end structure;

library IEEE;
use IEEE.std_logic_1164.all;

entity dff is
port(d, gclk, rnot: in STD_logic;
q: out STD_Logic);
end dff;
architecture structure of dff is
begin
start: process(gclk,rnot)
begin
if ( rising_edge(gclk) or rnot = '0') then
	if (rnot = '0') then
	q <= '0';
	else 
	q <= d;
	end if;
end if;
end process;
end structure;





library IEEE;

use IEEE.std_logic_1164.all;

package 
   CONV_PACK_top_g_hub_mux4_g_clock_freq200000000_g_color_depth8_g_num_row4_g_num_col4 
   is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type UNSIGNED is array (INTEGER range <>) of std_logic;
   
   -- Declarations for conversion functions.
   function BIT_to_std_logic(arg : in BIT) return std_logic;

end 
   CONV_PACK_top_g_hub_mux4_g_clock_freq200000000_g_color_depth8_g_num_row4_g_num_col4;

package body 
   CONV_PACK_top_g_hub_mux4_g_clock_freq200000000_g_color_depth8_g_num_row4_g_num_col4 
   is
   
   -- enum type to std_logic function
   function BIT_to_std_logic(arg : in BIT) return std_logic is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when '0' => return '0';
         when '1' => return '1';
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return '0';
      end case;
   end;

end 
   CONV_PACK_top_g_hub_mux4_g_clock_freq200000000_g_color_depth8_g_num_row4_g_num_col4;

library IEEE;

use IEEE.std_logic_1164.all;

use 
   work.CONV_PACK_top_g_hub_mux4_g_clock_freq200000000_g_color_depth8_g_num_row4_g_num_col4.all;

entity 
   top_g_hub_mux4_g_clock_freq200000000_g_color_depth8_g_num_row4_g_num_col4 is

   port( clk : in std_logic;  reset : in BIT;  top_data : in std_logic_vector 
         (23 downto 0);  top_dv_i, top_u_l : in std_logic;  top_ack : out 
         std_logic;  hub_mux_o : out UNSIGNED (3 downto 0);  hub_clk_o, 
         hub_latch_o, hub_blank_o, hub_g0_o, hub_b0_o, hub_r0_o : out std_logic
         );

end top_g_hub_mux4_g_clock_freq200000000_g_color_depth8_g_num_row4_g_num_col4;

architecture SYN_rtl of 
   top_g_hub_mux4_g_clock_freq200000000_g_color_depth8_g_num_row4_g_num_col4 is

   component inv
      port( inb : in std_logic;  outb : out std_logic);
   end component;
   
   component nor3
      port( a, b, c : in std_logic;  outb : out std_logic);
   end component;
   
   component nand2
      port( a, b : in std_logic;  outb : out std_logic);
   end component;
   
   component oai12
      port( b, c, a : in std_logic;  outb : out std_logic);
   end component;
   
   component nand3
      port( a, b, c : in std_logic;  outb : out std_logic);
   end component;
   
   component nand4
      port( a, b, c, d : in std_logic;  outb : out std_logic);
   end component;
   
   component nor2
      port( a, b : in std_logic;  outb : out std_logic);
   end component;
   
   component aoi22
      port( a, b, c, d : in std_logic;  outb : out std_logic);
   end component;
   
   component oai22
      port( a, b, c, d : in std_logic;  outb : out std_logic);
   end component;
   
   component aoi12
      port( b, c, a : in std_logic;  outb : out std_logic);
   end component;
   
   component xor2
      port( a, b : in std_logic;  outb : out std_logic);
   end component;
   
   component dff
      port( d, gclk, rnot : in std_logic;  q : out std_logic);
   end component;
   
   signal reset_port, top_ack_port, hub_mux_o_3_port, hub_mux_o_2_port, 
      hub_mux_o_1_port, hub_mux_o_0_port, hub_clk_o_port, hub_latch_o_port, 
      hub_blank_o_port, hub_g0_o_port, hub_b0_o_port, hub_r0_o_port, 
      mem_sipo_r0_7_port, mem_sipo_r0_6_port, mem_sipo_r0_5_port, 
      mem_sipo_r0_4_port, mem_sipo_r0_3_port, mem_sipo_r0_2_port, 
      mem_sipo_r0_1_port, mem_sipo_r0_0_port, mem_sipo_g0_7_port, 
      mem_sipo_g0_6_port, mem_sipo_g0_5_port, mem_sipo_g0_4_port, 
      mem_sipo_g0_3_port, mem_sipo_g0_2_port, mem_sipo_g0_1_port, 
      mem_sipo_g0_0_port, mem_sipo_b0_7_port, mem_sipo_b0_6_port, 
      mem_sipo_b0_5_port, mem_sipo_b0_4_port, mem_sipo_b0_3_port, 
      mem_sipo_b0_2_port, mem_sipo_b0_1_port, mem_sipo_b0_0_port, 
      mem_out_r0_7_port, mem_out_r0_6_port, mem_out_r0_5_port, 
      mem_out_r0_4_port, mem_out_r0_3_port, mem_out_r0_2_port, 
      mem_out_r0_1_port, mem_out_r0_0_port, mem_out_g0_7_port, 
      mem_out_g0_6_port, mem_out_g0_5_port, mem_out_g0_4_port, 
      mem_out_g0_3_port, mem_out_g0_2_port, mem_out_g0_1_port, 
      mem_out_g0_0_port, mem_out_b0_7_port, mem_out_b0_6_port, 
      mem_out_b0_5_port, mem_out_b0_4_port, mem_out_b0_3_port, 
      mem_out_b0_2_port, mem_out_b0_1_port, mem_out_b0_0_port, addr_i_3_port, 
      addr_i_2_port, addr_i_1_port, addr_i_0_port, reg_hub_f, hub_reg_f, 
      mem_reg_f, mem_hub_f, registers_n286, registers_n285, registers_n284, 
      registers_n283, registers_n282, registers_n281, registers_n280, 
      registers_n279, registers_n278, registers_n277, registers_n276, 
      registers_n275, registers_n274, registers_n273, registers_n272, 
      registers_n271, registers_n270, registers_n269, registers_n268, 
      registers_n267, registers_n266, registers_n265, registers_n264, 
      registers_n263, registers_n262, registers_n261, registers_n260, 
      registers_n259, registers_n258, registers_n257, registers_n256, 
      registers_n255, registers_n254, registers_n253, registers_n252, 
      registers_n251, registers_n250, registers_n249, registers_n248, 
      registers_n247, registers_n246, registers_n245, registers_n244, 
      registers_n243, registers_n242, registers_n241, registers_n240, 
      registers_n239, registers_n238, registers_n237, registers_n236, 
      registers_n235, registers_n234, registers_n233, registers_n232, 
      registers_n231, registers_n230, registers_n229, registers_n228, 
      registers_n227, registers_n226, registers_n225, registers_n224, 
      registers_n82, registers_n81, registers_n80, registers_n79, registers_n78
      , registers_n77, registers_n76, registers_n75, registers_n74, 
      registers_n73, registers_n72, registers_n71, registers_n70, registers_n69
      , registers_n68, registers_n67, registers_n66, registers_n65, 
      registers_n64, registers_n63, registers_n62, registers_n61, registers_n60
      , registers_n59, registers_n58, registers_n57, registers_n56, 
      registers_n55, registers_n54, registers_n53, registers_n52, registers_n51
      , registers_n50, registers_n49, registers_n48, registers_n47, 
      registers_n46, registers_n45, registers_n44, registers_n43, registers_n42
      , registers_n41, registers_n40, registers_n39, registers_n38, 
      registers_n37, registers_n36, registers_n35, registers_n34, registers_n33
      , registers_n32, registers_n31, registers_n30, registers_n29, 
      registers_n28, registers_n27, registers_n26, registers_n25, registers_n24
      , registers_n23, registers_n22, registers_n21, registers_n20, 
      registers_n19, registers_s_delay_0_port, registers_s_delay_1_port, 
      registers_s_mem_sipo_b0_0_port, registers_s_mem_sipo_b0_1_port, 
      registers_s_mem_sipo_b0_2_port, registers_s_mem_sipo_b0_3_port, 
      registers_s_mem_sipo_b0_4_port, registers_s_mem_sipo_b0_5_port, 
      registers_s_mem_sipo_b0_6_port, registers_s_mem_sipo_b0_7_port, 
      registers_s_mem_sipo_g0_0_port, registers_s_mem_sipo_g0_1_port, 
      registers_s_mem_sipo_g0_2_port, registers_s_mem_sipo_g0_3_port, 
      registers_s_mem_sipo_g0_4_port, registers_s_mem_sipo_g0_5_port, 
      registers_s_mem_sipo_g0_6_port, registers_s_mem_sipo_g0_7_port, 
      registers_s_mem_sipo_r0_0_port, registers_s_mem_sipo_r0_1_port, 
      registers_s_mem_sipo_r0_2_port, registers_s_mem_sipo_r0_3_port, 
      registers_s_mem_sipo_r0_4_port, registers_s_mem_sipo_r0_5_port, 
      registers_s_mem_sipo_r0_6_port, registers_s_mem_sipo_r0_7_port, 
      registers_reg_col_inc_0_port, registers_reg_col_inc_1_port, 
      registers_reg_cd_0_port, registers_reg_cd_1_port, registers_reg_cd_2_port
      , registers_reg_row_0_port, registers_reg_row_1_port, 
      registers_mem_to_reg_0_port, registers_mem_to_reg_1_port, 
      load_n_store_n303, load_n_store_n302, load_n_store_n301, 
      load_n_store_n300, load_n_store_n299, load_n_store_n92, load_n_store_n91,
      load_n_store_n90, load_n_store_n89, load_n_store_n88, load_n_store_n87, 
      load_n_store_n86, load_n_store_n85, load_n_store_n84, load_n_store_n83, 
      load_n_store_n82, load_n_store_n81, load_n_store_n80, load_n_store_n79, 
      load_n_store_n78, load_n_store_n77, load_n_store_n76, load_n_store_n75, 
      load_n_store_n74, load_n_store_n73, load_n_store_n72, load_n_store_n71, 
      load_n_store_n70, load_n_store_n69, load_n_store_n68, load_n_store_n67, 
      load_n_store_n66, load_n_store_n65, load_n_store_n64, load_n_store_n63, 
      load_n_store_n62, load_n_store_n61, load_n_store_n60, load_n_store_n59, 
      load_n_store_n58, load_n_store_n57, load_n_store_n56, load_n_store_n55, 
      load_n_store_n54, load_n_store_n53, load_n_store_n52, load_n_store_n51, 
      load_n_store_n50, load_n_store_n49, load_n_store_n48, load_n_store_n47, 
      load_n_store_n46, load_n_store_n45, load_n_store_n44, load_n_store_n43, 
      load_n_store_n42, load_n_store_n41, load_n_store_n40, load_n_store_n39, 
      load_n_store_n38, load_n_store_n37, load_n_store_n36, load_n_store_n35, 
      load_n_store_n34, load_n_store_n33, load_n_store_n32, load_n_store_n31, 
      load_n_store_n30, load_n_store_n29, load_n_store_n28, load_n_store_n27, 
      load_n_store_n26, load_n_store_n25, load_n_store_n24, load_n_store_n23, 
      load_n_store_n22, load_n_store_n21, load_n_store_n20, load_n_store_n19, 
      load_n_store_n18, load_n_store_n17, load_n_store_n16, load_n_store_n15, 
      load_n_store_n14, load_n_store_n13, load_n_store_n12, load_n_store_n11, 
      load_n_store_n10, load_n_store_n9, load_n_store_n8, load_n_store_n7, 
      load_n_store_mem_timer_0_port, load_n_store_mem_timer_1_port, 
      load_n_store_mem_timer_2_port, load_n_store_mem_timer_3_port, 
      load_n_store_mem_timer_4_port, load_n_store_mem_timer_5_port, 
      load_n_store_mem_timer_6_port, load_n_store_mem_timer_7_port, 
      load_n_store_mem_timer_8_port, load_n_store_mem_timer_9_port, 
      load_n_store_mem_timer_10_port, load_n_store_mem_timer_11_port, 
      load_n_store_mem_timer_12_port, load_n_store_mem_timer_13_port, 
      load_n_store_mem_timer_14_port, load_n_store_mem_timer_15_port, 
      load_n_store_mem_timer_16_port, load_n_store_mem_timer_17_port, 
      load_n_store_mem_timer_18_port, load_n_store_mem_timer_19_port, 
      load_n_store_mem_timer_20_port, load_n_store_mem_timer_21_port, 
      load_n_store_mem_timer_22_port, load_n_store_mem_timer_23_port, 
      load_n_store_mem_timer_24_port, load_n_store_mem_timer_25_port, 
      load_n_store_mem_timer_26_port, load_n_store_mem_timer_27_port, 
      load_n_store_mem_timer_28_port, load_n_store_mem_timer_29_port, 
      load_n_store_mem_timer_30_port, load_n_store_mem_timer_31_port, 
      load_n_store_simple_mem_sm_0_port, load_n_store_simple_mem_sm_1_port, 
      load_n_store_lazy_in_2_0_port, load_n_store_lazy_in_2_1_port, 
      load_n_store_lazy_in_2_2_port, load_n_store_lazy_in_2_3_port, 
      load_n_store_lazy_in_2_4_port, load_n_store_lazy_in_2_5_port, 
      load_n_store_lazy_in_2_6_port, load_n_store_lazy_in_2_7_port, 
      load_n_store_lazy_in_1_0_port, load_n_store_lazy_in_1_1_port, 
      load_n_store_lazy_in_1_2_port, load_n_store_lazy_in_1_3_port, 
      load_n_store_lazy_in_1_4_port, load_n_store_lazy_in_1_5_port, 
      load_n_store_lazy_in_1_6_port, load_n_store_lazy_in_1_7_port, 
      load_n_store_lazy_in_0_0_port, load_n_store_lazy_in_0_1_port, 
      load_n_store_lazy_in_0_2_port, load_n_store_lazy_in_0_3_port, 
      load_n_store_lazy_in_0_4_port, load_n_store_lazy_in_0_5_port, 
      load_n_store_lazy_in_0_6_port, load_n_store_lazy_in_0_7_port, 
      load_n_store_lazy_out_2_0_port, load_n_store_lazy_out_2_1_port, 
      load_n_store_lazy_out_2_2_port, load_n_store_lazy_out_2_3_port, 
      load_n_store_lazy_out_2_4_port, load_n_store_lazy_out_2_5_port, 
      load_n_store_lazy_out_2_6_port, load_n_store_lazy_out_2_7_port, 
      load_n_store_lazy_out_1_0_port, load_n_store_lazy_out_1_1_port, 
      load_n_store_lazy_out_1_2_port, load_n_store_lazy_out_1_3_port, 
      load_n_store_lazy_out_1_4_port, load_n_store_lazy_out_1_5_port, 
      load_n_store_lazy_out_1_6_port, load_n_store_lazy_out_1_7_port, 
      load_n_store_lazy_out_0_0_port, load_n_store_lazy_out_0_1_port, 
      load_n_store_lazy_out_0_2_port, load_n_store_lazy_out_0_3_port, 
      load_n_store_lazy_out_0_4_port, load_n_store_lazy_out_0_5_port, 
      load_n_store_lazy_out_0_6_port, load_n_store_lazy_out_0_7_port, 
      load_n_store_we_i, display_out_n912, display_out_n911, display_out_n910, 
      display_out_n909, display_out_n908, display_out_n907, display_out_n906, 
      display_out_n905, display_out_n904, display_out_n903, display_out_n902, 
      display_out_n901, display_out_n900, display_out_n899, display_out_n898, 
      display_out_n897, display_out_n896, display_out_n895, display_out_n894, 
      display_out_n893, display_out_n892, display_out_n891, display_out_n890, 
      display_out_n889, display_out_n888, display_out_n887, display_out_n886, 
      display_out_n885, display_out_n884, display_out_n883, display_out_n882, 
      display_out_n881, display_out_n880, display_out_n879, display_out_n878, 
      display_out_n877, display_out_n876, display_out_n875, display_out_n874, 
      display_out_n873, display_out_n872, display_out_n871, display_out_n870, 
      display_out_n869, display_out_n868, display_out_n867, display_out_n866, 
      display_out_n865, display_out_n864, display_out_n863, display_out_n862, 
      display_out_n861, display_out_n860, display_out_n859, display_out_n858, 
      display_out_n857, display_out_n856, display_out_n855, display_out_n854, 
      display_out_n853, display_out_n852, display_out_n851, display_out_n850, 
      display_out_n849, display_out_n848, display_out_n847, display_out_n846, 
      display_out_n845, display_out_n844, display_out_n843, display_out_n842, 
      display_out_n841, display_out_n840, display_out_n839, display_out_n838, 
      display_out_n837, display_out_n836, display_out_n835, display_out_n834, 
      display_out_n833, display_out_n832, display_out_n831, display_out_n830, 
      display_out_n829, display_out_n828, display_out_n827, display_out_n826, 
      display_out_n825, display_out_n824, display_out_n823, display_out_n822, 
      display_out_n821, display_out_n820, display_out_n819, display_out_n818, 
      display_out_n817, display_out_n816, display_out_n815, display_out_n814, 
      display_out_n813, display_out_n812, display_out_n811, display_out_n810, 
      display_out_n809, display_out_n808, display_out_n807, display_out_n806, 
      display_out_n805, display_out_n804, display_out_n803, display_out_n802, 
      display_out_n801, display_out_n800, display_out_n799, display_out_n798, 
      display_out_n797, display_out_n256, display_out_n255, display_out_n254, 
      display_out_n253, display_out_n252, display_out_n251, display_out_n250, 
      display_out_n249, display_out_n248, display_out_n247, display_out_n246, 
      display_out_n245, display_out_n244, display_out_n243, display_out_n242, 
      display_out_n241, display_out_n240, display_out_n239, display_out_n238, 
      display_out_n237, display_out_n236, display_out_n235, display_out_n234, 
      display_out_n233, display_out_n232, display_out_n231, display_out_n230, 
      display_out_n229, display_out_n228, display_out_n227, display_out_n226, 
      display_out_n225, display_out_n224, display_out_n223, display_out_n222, 
      display_out_n221, display_out_n220, display_out_n219, display_out_n218, 
      display_out_n217, display_out_n216, display_out_n215, display_out_n214, 
      display_out_n213, display_out_n212, display_out_n211, display_out_n210, 
      display_out_n209, display_out_n208, display_out_n207, display_out_n206, 
      display_out_n205, display_out_n204, display_out_n203, display_out_n202, 
      display_out_n201, display_out_n200, display_out_n199, display_out_n198, 
      display_out_n197, display_out_n196, display_out_n195, display_out_n194, 
      display_out_n193, display_out_n192, display_out_n191, display_out_n190, 
      display_out_n189, display_out_n188, display_out_n187, display_out_n186, 
      display_out_n185, display_out_n184, display_out_n183, display_out_n182, 
      display_out_n181, display_out_n180, display_out_n179, display_out_n178, 
      display_out_n177, display_out_n176, display_out_n175, display_out_n174, 
      display_out_n173, display_out_n172, display_out_n171, display_out_n170, 
      display_out_n169, display_out_n168, display_out_n167, display_out_n166, 
      display_out_n165, display_out_n164, display_out_n163, display_out_n162, 
      display_out_n161, display_out_n160, display_out_n159, display_out_n158, 
      display_out_n157, display_out_n156, display_out_n155, display_out_n154, 
      display_out_n153, display_out_n152, display_out_n151, display_out_n150, 
      display_out_n149, display_out_n148, display_out_n147, display_out_n146, 
      display_out_n145, display_out_n144, display_out_n143, display_out_n142, 
      display_out_n141, display_out_n140, display_out_n139, display_out_n138, 
      display_out_n137, display_out_n136, display_out_n135, display_out_n134, 
      display_out_n133, display_out_n132, display_out_n131, display_out_n130, 
      display_out_n129, display_out_n128, display_out_n127, display_out_n126, 
      display_out_n125, display_out_n124, display_out_n123, display_out_n122, 
      display_out_n121, display_out_n120, display_out_n119, display_out_n118, 
      display_out_n117, display_out_n116, display_out_n115, display_out_n114, 
      display_out_n113, display_out_n112, display_out_n111, display_out_n110, 
      display_out_n109, display_out_n108, display_out_n107, display_out_n106, 
      display_out_n105, display_out_n104, display_out_n103, display_out_n102, 
      display_out_n101, display_out_n100, display_out_n99, display_out_n98, 
      display_out_n97, display_out_n96, display_out_n95, display_out_n94, 
      display_out_n93, display_out_n92, display_out_n91, display_out_n90, 
      display_out_n89, display_out_n88, display_out_hub_piso_b0_0_port, 
      display_out_hub_piso_b0_1_port, display_out_hub_piso_b0_2_port, 
      display_out_hub_piso_b0_3_port, display_out_hub_piso_b0_4_port, 
      display_out_hub_piso_b0_5_port, display_out_hub_piso_b0_6_port, 
      display_out_hub_piso_b0_7_port, display_out_hub_piso_g0_0_port, 
      display_out_hub_piso_g0_1_port, display_out_hub_piso_g0_2_port, 
      display_out_hub_piso_g0_3_port, display_out_hub_piso_g0_4_port, 
      display_out_hub_piso_g0_5_port, display_out_hub_piso_g0_6_port, 
      display_out_hub_piso_g0_7_port, display_out_hub_piso_r0_0_port, 
      display_out_hub_piso_r0_1_port, display_out_hub_piso_r0_2_port, 
      display_out_hub_piso_r0_3_port, display_out_hub_piso_r0_4_port, 
      display_out_hub_piso_r0_5_port, display_out_hub_piso_r0_6_port, 
      display_out_hub_piso_r0_7_port, display_out_clk_timer_0_port, 
      display_out_clk_timer_1_port, display_out_clk_timer_2_port, 
      display_out_clk_timer_3_port, display_out_clk_timer_4_port, 
      display_out_clk_timer_5_port, display_out_clk_timer_6_port, 
      display_out_clk_timer_7_port, display_out_clk_timer_8_port, 
      display_out_clk_timer_9_port, display_out_clk_timer_10_port, 
      display_out_clk_timer_11_port, display_out_clk_timer_12_port, 
      display_out_clk_timer_13_port, display_out_clk_timer_14_port, 
      display_out_clk_timer_15_port, display_out_clk_timer_16_port, 
      display_out_clk_timer_17_port, display_out_clk_timer_18_port, 
      display_out_clk_timer_19_port, display_out_clk_timer_20_port, 
      display_out_clk_timer_21_port, display_out_clk_timer_22_port, 
      display_out_clk_timer_23_port, display_out_clk_timer_24_port, 
      display_out_clk_timer_25_port, display_out_clk_timer_26_port, 
      display_out_clk_timer_27_port, display_out_clk_timer_28_port, 
      display_out_clk_timer_29_port, display_out_clk_timer_30_port, 
      display_out_clk_timer_31_port, display_out_disp_timer_0_port, 
      display_out_disp_timer_1_port, display_out_disp_timer_2_port, 
      display_out_disp_timer_3_port, display_out_disp_timer_4_port, 
      display_out_disp_timer_5_port, display_out_disp_timer_6_port, 
      display_out_disp_timer_7_port, display_out_disp_timer_8_port, 
      display_out_disp_timer_9_port, display_out_disp_timer_10_port, 
      display_out_disp_timer_11_port, display_out_disp_timer_12_port, 
      display_out_disp_timer_13_port, display_out_disp_timer_14_port, 
      display_out_disp_timer_15_port, display_out_disp_timer_16_port, 
      display_out_disp_timer_17_port, display_out_disp_timer_18_port, 
      display_out_disp_timer_19_port, display_out_disp_timer_20_port, 
      display_out_disp_timer_21_port, display_out_disp_timer_22_port, 
      display_out_disp_timer_23_port, display_out_disp_timer_24_port, 
      display_out_disp_timer_25_port, display_out_disp_timer_26_port, 
      display_out_disp_timer_27_port, display_out_disp_timer_28_port, 
      display_out_disp_timer_29_port, display_out_disp_timer_30_port, 
      display_out_disp_timer_31_port, display_out_h_col_0_port, 
      display_out_h_col_1_port, display_out_h_col_2_port, 
      display_out_h_col_3_port, display_out_h_col_4_port, 
      display_out_h_col_5_port, display_out_h_col_6_port, 
      display_out_h_col_7_port, display_out_h_col_8_port, 
      display_out_h_col_9_port, display_out_h_col_10_port, 
      display_out_h_col_11_port, display_out_h_col_12_port, 
      display_out_h_col_13_port, display_out_h_col_14_port, 
      display_out_h_col_15_port, display_out_h_col_16_port, 
      display_out_h_col_17_port, display_out_h_col_18_port, 
      display_out_h_col_19_port, display_out_h_col_20_port, 
      display_out_h_col_21_port, display_out_h_col_22_port, 
      display_out_h_col_23_port, display_out_h_col_24_port, 
      display_out_h_col_25_port, display_out_h_col_26_port, 
      display_out_h_col_27_port, display_out_h_col_28_port, 
      display_out_h_col_29_port, display_out_h_col_30_port, 
      display_out_h_col_31_port, display_out_h_row_0_port, 
      display_out_h_row_1_port, display_out_h_row_2_port, 
      display_out_h_row_3_port, display_out_h_row_4_port, 
      display_out_h_row_5_port, display_out_h_row_6_port, 
      display_out_h_row_7_port, display_out_h_row_8_port, 
      display_out_h_row_9_port, display_out_h_row_10_port, 
      display_out_h_row_11_port, display_out_h_row_12_port, 
      display_out_h_row_13_port, display_out_h_row_14_port, 
      display_out_h_row_15_port, display_out_h_row_16_port, 
      display_out_h_row_17_port, display_out_h_row_18_port, 
      display_out_h_row_19_port, display_out_h_row_20_port, 
      display_out_h_row_21_port, display_out_h_row_22_port, 
      display_out_h_row_23_port, display_out_h_row_24_port, 
      display_out_h_row_25_port, display_out_h_row_26_port, 
      display_out_h_row_27_port, display_out_h_row_28_port, 
      display_out_h_row_29_port, display_out_h_row_30_port, 
      display_out_h_row_31_port, display_out_bcd_time_0_port, 
      display_out_bcd_time_1_port, display_out_bcd_time_2_port, 
      display_out_hub_out_sm_0_port, display_out_hub_out_sm_1_port, 
      display_out_hub_out_sm_2_port, load_n_store_RGB_Array_0_n600, 
      load_n_store_RGB_Array_0_n599, load_n_store_RGB_Array_0_n598, 
      load_n_store_RGB_Array_0_n597, load_n_store_RGB_Array_0_n596, 
      load_n_store_RGB_Array_0_n595, load_n_store_RGB_Array_0_n594, 
      load_n_store_RGB_Array_0_n593, load_n_store_RGB_Array_0_n592, 
      load_n_store_RGB_Array_0_n591, load_n_store_RGB_Array_0_n590, 
      load_n_store_RGB_Array_0_n589, load_n_store_RGB_Array_0_n588, 
      load_n_store_RGB_Array_0_n587, load_n_store_RGB_Array_0_n586, 
      load_n_store_RGB_Array_0_n585, load_n_store_RGB_Array_0_n584, 
      load_n_store_RGB_Array_0_n583, load_n_store_RGB_Array_0_n582, 
      load_n_store_RGB_Array_0_n581, load_n_store_RGB_Array_0_n580, 
      load_n_store_RGB_Array_0_n579, load_n_store_RGB_Array_0_n578, 
      load_n_store_RGB_Array_0_n577, load_n_store_RGB_Array_0_n576, 
      load_n_store_RGB_Array_0_n575, load_n_store_RGB_Array_0_n574, 
      load_n_store_RGB_Array_0_n573, load_n_store_RGB_Array_0_n572, 
      load_n_store_RGB_Array_0_n571, load_n_store_RGB_Array_0_n570, 
      load_n_store_RGB_Array_0_n569, load_n_store_RGB_Array_0_n568, 
      load_n_store_RGB_Array_0_n567, load_n_store_RGB_Array_0_n566, 
      load_n_store_RGB_Array_0_n565, load_n_store_RGB_Array_0_n564, 
      load_n_store_RGB_Array_0_n563, load_n_store_RGB_Array_0_n562, 
      load_n_store_RGB_Array_0_n561, load_n_store_RGB_Array_0_n560, 
      load_n_store_RGB_Array_0_n559, load_n_store_RGB_Array_0_n558, 
      load_n_store_RGB_Array_0_n557, load_n_store_RGB_Array_0_n556, 
      load_n_store_RGB_Array_0_n555, load_n_store_RGB_Array_0_n554, 
      load_n_store_RGB_Array_0_n553, load_n_store_RGB_Array_0_n552, 
      load_n_store_RGB_Array_0_n551, load_n_store_RGB_Array_0_n550, 
      load_n_store_RGB_Array_0_n549, load_n_store_RGB_Array_0_n548, 
      load_n_store_RGB_Array_0_n547, load_n_store_RGB_Array_0_n546, 
      load_n_store_RGB_Array_0_n545, load_n_store_RGB_Array_0_n544, 
      load_n_store_RGB_Array_0_n543, load_n_store_RGB_Array_0_n542, 
      load_n_store_RGB_Array_0_n541, load_n_store_RGB_Array_0_n540, 
      load_n_store_RGB_Array_0_n539, load_n_store_RGB_Array_0_n538, 
      load_n_store_RGB_Array_0_n537, load_n_store_RGB_Array_0_n536, 
      load_n_store_RGB_Array_0_n535, load_n_store_RGB_Array_0_n534, 
      load_n_store_RGB_Array_0_n533, load_n_store_RGB_Array_0_n532, 
      load_n_store_RGB_Array_0_n531, load_n_store_RGB_Array_0_n530, 
      load_n_store_RGB_Array_0_n529, load_n_store_RGB_Array_0_n528, 
      load_n_store_RGB_Array_0_n527, load_n_store_RGB_Array_0_n526, 
      load_n_store_RGB_Array_0_n525, load_n_store_RGB_Array_0_n524, 
      load_n_store_RGB_Array_0_n523, load_n_store_RGB_Array_0_n522, 
      load_n_store_RGB_Array_0_n521, load_n_store_RGB_Array_0_n520, 
      load_n_store_RGB_Array_0_n519, load_n_store_RGB_Array_0_n518, 
      load_n_store_RGB_Array_0_n517, load_n_store_RGB_Array_0_n516, 
      load_n_store_RGB_Array_0_n515, load_n_store_RGB_Array_0_n514, 
      load_n_store_RGB_Array_0_n513, load_n_store_RGB_Array_0_n512, 
      load_n_store_RGB_Array_0_n511, load_n_store_RGB_Array_0_n510, 
      load_n_store_RGB_Array_0_n509, load_n_store_RGB_Array_0_n508, 
      load_n_store_RGB_Array_0_n507, load_n_store_RGB_Array_0_n506, 
      load_n_store_RGB_Array_0_n505, load_n_store_RGB_Array_0_n504, 
      load_n_store_RGB_Array_0_n503, load_n_store_RGB_Array_0_n502, 
      load_n_store_RGB_Array_0_n501, load_n_store_RGB_Array_0_n500, 
      load_n_store_RGB_Array_0_n499, load_n_store_RGB_Array_0_n498, 
      load_n_store_RGB_Array_0_n497, load_n_store_RGB_Array_0_n496, 
      load_n_store_RGB_Array_0_n495, load_n_store_RGB_Array_0_n494, 
      load_n_store_RGB_Array_0_n493, load_n_store_RGB_Array_0_n492, 
      load_n_store_RGB_Array_0_n491, load_n_store_RGB_Array_0_n490, 
      load_n_store_RGB_Array_0_n489, load_n_store_RGB_Array_0_n488, 
      load_n_store_RGB_Array_0_n487, load_n_store_RGB_Array_0_n486, 
      load_n_store_RGB_Array_0_n485, load_n_store_RGB_Array_0_n484, 
      load_n_store_RGB_Array_0_n483, load_n_store_RGB_Array_0_n482, 
      load_n_store_RGB_Array_0_n481, load_n_store_RGB_Array_0_n480, 
      load_n_store_RGB_Array_0_n479, load_n_store_RGB_Array_0_n478, 
      load_n_store_RGB_Array_0_n477, load_n_store_RGB_Array_0_n476, 
      load_n_store_RGB_Array_0_n475, load_n_store_RGB_Array_0_n474, 
      load_n_store_RGB_Array_0_n473, load_n_store_RGB_Array_0_n472, 
      load_n_store_RGB_Array_0_n471, load_n_store_RGB_Array_0_n470, 
      load_n_store_RGB_Array_0_n469, load_n_store_RGB_Array_0_n468, 
      load_n_store_RGB_Array_0_n467, load_n_store_RGB_Array_0_n466, 
      load_n_store_RGB_Array_0_n465, load_n_store_RGB_Array_0_n464, 
      load_n_store_RGB_Array_0_n463, load_n_store_RGB_Array_0_n462, 
      load_n_store_RGB_Array_0_n461, load_n_store_RGB_Array_0_n460, 
      load_n_store_RGB_Array_0_n459, load_n_store_RGB_Array_0_n458, 
      load_n_store_RGB_Array_0_n457, load_n_store_RGB_Array_0_n456, 
      load_n_store_RGB_Array_0_n455, load_n_store_RGB_Array_0_n454, 
      load_n_store_RGB_Array_0_n453, load_n_store_RGB_Array_0_n452, 
      load_n_store_RGB_Array_0_n451, load_n_store_RGB_Array_0_n450, 
      load_n_store_RGB_Array_0_n449, load_n_store_RGB_Array_0_n448, 
      load_n_store_RGB_Array_0_n447, load_n_store_RGB_Array_0_n446, 
      load_n_store_RGB_Array_0_n445, load_n_store_RGB_Array_0_n444, 
      load_n_store_RGB_Array_0_n443, load_n_store_RGB_Array_0_n442, 
      load_n_store_RGB_Array_0_n441, load_n_store_RGB_Array_0_n440, 
      load_n_store_RGB_Array_0_n439, load_n_store_RGB_Array_0_n438, 
      load_n_store_RGB_Array_0_n437, load_n_store_RGB_Array_0_n436, 
      load_n_store_RGB_Array_0_n435, load_n_store_RGB_Array_0_n434, 
      load_n_store_RGB_Array_0_n433, load_n_store_RGB_Array_0_n432, 
      load_n_store_RGB_Array_0_n431, load_n_store_RGB_Array_0_n430, 
      load_n_store_RGB_Array_0_n429, load_n_store_RGB_Array_0_n428, 
      load_n_store_RGB_Array_0_n427, load_n_store_RGB_Array_0_n426, 
      load_n_store_RGB_Array_0_n425, load_n_store_RGB_Array_0_n424, 
      load_n_store_RGB_Array_0_n423, load_n_store_RGB_Array_0_n422, 
      load_n_store_RGB_Array_0_n421, load_n_store_RGB_Array_0_n420, 
      load_n_store_RGB_Array_0_n419, load_n_store_RGB_Array_0_n418, 
      load_n_store_RGB_Array_0_n417, load_n_store_RGB_Array_0_n416, 
      load_n_store_RGB_Array_0_n415, load_n_store_RGB_Array_0_n414, 
      load_n_store_RGB_Array_0_n413, load_n_store_RGB_Array_0_n412, 
      load_n_store_RGB_Array_0_n411, load_n_store_RGB_Array_0_n410, 
      load_n_store_RGB_Array_0_n409, load_n_store_RGB_Array_0_n408, 
      load_n_store_RGB_Array_0_n407, load_n_store_RGB_Array_0_n406, 
      load_n_store_RGB_Array_0_n405, load_n_store_RGB_Array_0_n404, 
      load_n_store_RGB_Array_0_n403, load_n_store_RGB_Array_0_n402, 
      load_n_store_RGB_Array_0_n401, load_n_store_RGB_Array_0_n400, 
      load_n_store_RGB_Array_0_n399, load_n_store_RGB_Array_0_n398, 
      load_n_store_RGB_Array_0_n397, load_n_store_RGB_Array_0_n396, 
      load_n_store_RGB_Array_0_n395, load_n_store_RGB_Array_0_n394, 
      load_n_store_RGB_Array_0_n393, load_n_store_RGB_Array_0_n392, 
      load_n_store_RGB_Array_0_n391, load_n_store_RGB_Array_0_n390, 
      load_n_store_RGB_Array_0_n389, load_n_store_RGB_Array_0_n388, 
      load_n_store_RGB_Array_0_n387, load_n_store_RGB_Array_0_n386, 
      load_n_store_RGB_Array_0_n385, load_n_store_RGB_Array_0_n384, 
      load_n_store_RGB_Array_0_n383, load_n_store_RGB_Array_0_n382, 
      load_n_store_RGB_Array_0_n381, load_n_store_RGB_Array_0_n380, 
      load_n_store_RGB_Array_0_n379, load_n_store_RGB_Array_0_n378, 
      load_n_store_RGB_Array_0_n377, load_n_store_RGB_Array_0_n376, 
      load_n_store_RGB_Array_0_n375, load_n_store_RGB_Array_0_n374, 
      load_n_store_RGB_Array_0_n373, load_n_store_RGB_Array_0_n372, 
      load_n_store_RGB_Array_0_n371, load_n_store_RGB_Array_0_n370, 
      load_n_store_RGB_Array_0_n369, load_n_store_RGB_Array_0_n368, 
      load_n_store_RGB_Array_0_n367, load_n_store_RGB_Array_0_n366, 
      load_n_store_RGB_Array_0_n365, load_n_store_RGB_Array_0_n364, 
      load_n_store_RGB_Array_0_n363, load_n_store_RGB_Array_0_n362, 
      load_n_store_RGB_Array_0_n361, load_n_store_RGB_Array_0_n360, 
      load_n_store_RGB_Array_0_n359, load_n_store_RGB_Array_0_n358, 
      load_n_store_RGB_Array_0_n357, load_n_store_RGB_Array_0_n356, 
      load_n_store_RGB_Array_0_n355, load_n_store_RGB_Array_0_n354, 
      load_n_store_RGB_Array_0_n353, load_n_store_RGB_Array_0_n352, 
      load_n_store_RGB_Array_0_n350, load_n_store_RGB_Array_0_n349, 
      load_n_store_RGB_Array_0_n347, load_n_store_RGB_Array_0_n346, 
      load_n_store_RGB_Array_0_n344, load_n_store_RGB_Array_0_n343, 
      load_n_store_RGB_Array_0_n341, load_n_store_RGB_Array_0_n340, 
      load_n_store_RGB_Array_0_n338, load_n_store_RGB_Array_0_n337, 
      load_n_store_RGB_Array_0_n335, load_n_store_RGB_Array_0_n334, 
      load_n_store_RGB_Array_0_n332, load_n_store_RGB_Array_0_n331, 
      load_n_store_RGB_Array_0_n329, load_n_store_RGB_Array_0_n174, 
      load_n_store_RGB_Array_0_n151, load_n_store_RGB_Array_0_n128, 
      load_n_store_RGB_Array_0_n105, load_n_store_RGB_Array_0_n82, 
      load_n_store_RGB_Array_0_n59, load_n_store_RGB_Array_0_n36, 
      load_n_store_RGB_Array_0_n2, 
      load_n_store_RGB_Array_0_block_ram_r_0_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_0_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_0_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_0_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_0_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_0_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_0_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_0_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_1_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_1_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_1_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_1_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_1_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_1_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_1_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_1_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_2_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_2_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_2_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_2_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_2_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_2_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_2_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_2_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_3_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_3_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_3_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_3_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_3_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_3_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_3_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_3_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_4_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_4_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_4_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_4_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_4_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_4_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_4_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_4_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_5_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_5_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_5_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_5_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_5_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_5_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_5_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_5_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_6_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_6_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_6_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_6_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_6_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_6_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_6_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_6_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_7_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_7_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_7_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_7_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_7_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_7_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_7_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_7_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_8_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_8_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_8_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_8_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_8_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_8_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_8_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_8_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_9_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_9_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_9_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_9_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_9_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_9_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_9_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_9_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_10_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_10_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_10_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_10_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_10_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_10_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_10_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_10_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_11_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_11_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_11_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_11_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_11_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_11_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_11_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_11_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_12_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_12_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_12_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_12_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_12_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_12_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_12_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_12_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_13_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_13_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_13_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_13_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_13_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_13_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_13_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_13_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_14_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_14_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_14_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_14_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_14_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_14_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_14_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_14_7_port, 
      load_n_store_RGB_Array_0_block_ram_r_15_0_port, 
      load_n_store_RGB_Array_0_block_ram_r_15_1_port, 
      load_n_store_RGB_Array_0_block_ram_r_15_2_port, 
      load_n_store_RGB_Array_0_block_ram_r_15_3_port, 
      load_n_store_RGB_Array_0_block_ram_r_15_4_port, 
      load_n_store_RGB_Array_0_block_ram_r_15_5_port, 
      load_n_store_RGB_Array_0_block_ram_r_15_6_port, 
      load_n_store_RGB_Array_0_block_ram_r_15_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_0_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_0_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_0_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_0_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_0_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_0_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_0_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_0_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_1_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_1_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_1_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_1_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_1_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_1_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_1_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_1_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_2_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_2_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_2_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_2_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_2_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_2_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_2_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_2_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_3_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_3_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_3_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_3_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_3_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_3_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_3_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_3_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_4_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_4_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_4_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_4_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_4_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_4_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_4_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_4_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_5_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_5_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_5_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_5_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_5_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_5_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_5_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_5_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_6_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_6_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_6_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_6_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_6_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_6_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_6_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_6_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_7_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_7_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_7_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_7_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_7_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_7_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_7_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_7_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_8_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_8_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_8_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_8_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_8_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_8_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_8_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_8_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_9_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_9_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_9_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_9_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_9_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_9_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_9_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_9_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_10_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_10_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_10_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_10_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_10_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_10_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_10_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_10_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_11_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_11_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_11_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_11_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_11_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_11_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_11_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_11_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_12_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_12_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_12_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_12_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_12_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_12_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_12_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_12_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_13_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_13_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_13_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_13_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_13_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_13_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_13_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_13_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_14_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_14_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_14_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_14_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_14_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_14_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_14_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_14_7_port, 
      load_n_store_RGB_Array_2_block_ram_r_15_0_port, 
      load_n_store_RGB_Array_2_block_ram_r_15_1_port, 
      load_n_store_RGB_Array_2_block_ram_r_15_2_port, 
      load_n_store_RGB_Array_2_block_ram_r_15_3_port, 
      load_n_store_RGB_Array_2_block_ram_r_15_4_port, 
      load_n_store_RGB_Array_2_block_ram_r_15_5_port, 
      load_n_store_RGB_Array_2_block_ram_r_15_6_port, 
      load_n_store_RGB_Array_2_block_ram_r_15_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_0_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_0_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_0_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_0_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_0_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_0_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_0_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_0_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_1_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_1_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_1_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_1_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_1_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_1_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_1_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_1_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_2_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_2_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_2_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_2_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_2_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_2_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_2_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_2_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_3_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_3_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_3_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_3_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_3_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_3_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_3_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_3_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_4_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_4_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_4_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_4_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_4_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_4_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_4_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_4_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_5_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_5_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_5_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_5_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_5_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_5_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_5_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_5_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_6_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_6_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_6_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_6_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_6_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_6_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_6_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_6_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_7_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_7_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_7_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_7_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_7_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_7_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_7_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_7_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_8_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_8_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_8_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_8_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_8_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_8_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_8_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_8_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_9_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_9_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_9_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_9_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_9_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_9_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_9_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_9_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_10_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_10_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_10_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_10_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_10_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_10_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_10_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_10_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_11_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_11_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_11_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_11_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_11_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_11_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_11_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_11_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_12_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_12_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_12_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_12_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_12_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_12_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_12_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_12_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_13_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_13_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_13_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_13_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_13_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_13_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_13_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_13_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_14_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_14_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_14_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_14_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_14_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_14_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_14_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_14_7_port, 
      load_n_store_RGB_Array_1_block_ram_r_15_0_port, 
      load_n_store_RGB_Array_1_block_ram_r_15_1_port, 
      load_n_store_RGB_Array_1_block_ram_r_15_2_port, 
      load_n_store_RGB_Array_1_block_ram_r_15_3_port, 
      load_n_store_RGB_Array_1_block_ram_r_15_4_port, 
      load_n_store_RGB_Array_1_block_ram_r_15_5_port, 
      load_n_store_RGB_Array_1_block_ram_r_15_6_port, 
      load_n_store_RGB_Array_1_block_ram_r_15_7_port, n1, n2, n3, n4, n5, n6, 
      n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
      n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
      n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, 
      n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
      n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, 
      n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, 
      n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, 
      n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, 
      n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, 
      n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, 
      n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, 
      n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, 
      n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, 
      n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, 
      n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, 
      n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, 
      n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, 
      n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, 
      n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, 
      n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, 
      n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, 
      n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, 
      n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, 
      n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, 
      n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, 
      n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, 
      n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, 
      n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, 
      n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, 
      n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, 
      n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, 
      n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, 
      n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, 
      n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, 
      n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, 
      n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, 
      n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, 
      n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, 
      n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, 
      n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, 
      n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, 
      n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, 
      n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, 
      n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, 
      n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, 
      n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, 
      n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, 
      n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, 
      n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, 
      n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, 
      n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, 
      n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, 
      n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, 
      n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, 
      n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, 
      n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, 
      n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, 
      n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, 
      n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, 
      n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, 
      n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, 
      n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, 
      n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, 
      n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, 
      n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, 
      n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, 
      n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, 
      n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, 
      n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, 
      n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, 
      n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, 
      n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, 
      n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, 
      n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, 
      n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, 
      n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, 
      n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, 
      n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, 
      n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, 
      n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
      n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, 
      n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, 
      n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, 
      n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, 
      n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, 
      n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
      n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
      n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
      n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
      n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, 
      n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
      n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, 
      n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, 
      n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
      n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
      n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
      n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
      n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
      n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
      n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
      n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
      n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, 
      n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
      n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
      n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, 
      n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, 
      n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, 
      n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, 
      n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, 
      n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, 
      n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, 
      n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, 
      n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, 
      n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, 
      n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, 
      n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, 
      n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, 
      n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, 
      n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, 
      n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, 
      n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, 
      n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, 
      n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, 
      n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, 
      n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, 
      n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, 
      n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
      n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, 
      n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, 
      n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, 
      n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, 
      n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, 
      n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, 
      n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, 
      n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, 
      n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, 
      n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, 
      n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, 
      n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, 
      n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, 
      n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, 
      n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, 
      n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, 
      n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, 
      n2567, n2568, n2569, n2570, n2571, n2572 : std_logic;

begin
   reset_port <= BIT_to_std_logic(reset);
   top_ack <= top_ack_port;
   hub_mux_o <= ( hub_mux_o_3_port, hub_mux_o_2_port, hub_mux_o_1_port, 
      hub_mux_o_0_port );
   hub_clk_o <= hub_clk_o_port;
   hub_latch_o <= hub_latch_o_port;
   hub_blank_o <= hub_blank_o_port;
   hub_g0_o <= hub_g0_o_port;
   hub_b0_o <= hub_b0_o_port;
   hub_r0_o <= hub_r0_o_port;
   
   registers_n82 <= '1';
   registers_n81 <= '1';
   registers_n80 <= '1';
   registers_n79 <= '1';
   registers_n78 <= '1';
   registers_n77 <= '1';
   registers_n76 <= '1';
   registers_n75 <= '1';
   registers_n74 <= '1';
   registers_n73 <= '1';
   registers_n72 <= '1';
   registers_n71 <= '1';
   registers_n70 <= '1';
   registers_n69 <= '1';
   registers_n68 <= '1';
   registers_n67 <= '1';
   registers_n66 <= '1';
   registers_n65 <= '1';
   registers_n64 <= '1';
   registers_n63 <= '1';
   registers_n62 <= '1';
   registers_n61 <= '1';
   registers_n60 <= '1';
   registers_n59 <= '1';
   registers_n58 <= '1';
   registers_n57 <= '1';
   registers_n56 <= '1';
   registers_n55 <= '1';
   registers_n54 <= '1';
   registers_n53 <= '1';
   registers_n52 <= '1';
   registers_n51 <= '1';
   registers_n50 <= '1';
   registers_n49 <= '1';
   registers_n48 <= '1';
   registers_n47 <= '1';
   registers_n46 <= '1';
   registers_n45 <= '1';
   registers_n44 <= '1';
   registers_n43 <= '1';
   registers_n42 <= '1';
   registers_n41 <= '1';
   registers_n40 <= '1';
   registers_n39 <= '1';
   registers_n38 <= '1';
   registers_n37 <= '1';
   registers_n36 <= '1';
   registers_n35 <= '1';
   registers_n34 <= '1';
   registers_n33 <= '1';
   registers_n32 <= '1';
   registers_n31 <= '1';
   registers_n30 <= '1';
   registers_n29 <= '1';
   registers_n28 <= '1';
   registers_n27 <= '1';
   registers_n26 <= '1';
   registers_n25 <= '1';
   registers_n24 <= '1';
   registers_n23 <= '1';
   registers_n22 <= '1';
   registers_n21 <= '1';
   registers_n20 <= '1';
   registers_n19 <= '1';
   registers_mem_sipo_g0_reg_0_inst : dff port map( d => registers_n224, gclk 
                           => clk, rnot => registers_n19, q => 
                           mem_sipo_g0_0_port);
   registers_mem_sipo_g0_reg_1_inst : dff port map( d => registers_n225, gclk 
                           => clk, rnot => registers_n20, q => 
                           mem_sipo_g0_1_port);
   registers_mem_sipo_g0_reg_2_inst : dff port map( d => registers_n226, gclk 
                           => clk, rnot => registers_n21, q => 
                           mem_sipo_g0_2_port);
   registers_mem_sipo_g0_reg_3_inst : dff port map( d => registers_n227, gclk 
                           => clk, rnot => registers_n22, q => 
                           mem_sipo_g0_3_port);
   registers_mem_sipo_g0_reg_4_inst : dff port map( d => registers_n228, gclk 
                           => clk, rnot => registers_n23, q => 
                           mem_sipo_g0_4_port);
   registers_mem_sipo_g0_reg_5_inst : dff port map( d => registers_n229, gclk 
                           => clk, rnot => registers_n24, q => 
                           mem_sipo_g0_5_port);
   registers_mem_sipo_g0_reg_6_inst : dff port map( d => registers_n230, gclk 
                           => clk, rnot => registers_n25, q => 
                           mem_sipo_g0_6_port);
   registers_mem_sipo_g0_reg_7_inst : dff port map( d => registers_n231, gclk 
                           => clk, rnot => registers_n26, q => 
                           mem_sipo_g0_7_port);
   registers_mem_sipo_r0_reg_0_inst : dff port map( d => registers_n232, gclk 
                           => clk, rnot => registers_n27, q => 
                           mem_sipo_r0_0_port);
   registers_mem_sipo_r0_reg_1_inst : dff port map( d => registers_n233, gclk 
                           => clk, rnot => registers_n28, q => 
                           mem_sipo_r0_1_port);
   registers_mem_sipo_r0_reg_2_inst : dff port map( d => registers_n234, gclk 
                           => clk, rnot => registers_n29, q => 
                           mem_sipo_r0_2_port);
   registers_mem_sipo_r0_reg_3_inst : dff port map( d => registers_n235, gclk 
                           => clk, rnot => registers_n30, q => 
                           mem_sipo_r0_3_port);
   registers_mem_sipo_r0_reg_4_inst : dff port map( d => registers_n236, gclk 
                           => clk, rnot => registers_n31, q => 
                           mem_sipo_r0_4_port);
   registers_mem_sipo_r0_reg_5_inst : dff port map( d => registers_n237, gclk 
                           => clk, rnot => registers_n32, q => 
                           mem_sipo_r0_5_port);
   registers_mem_sipo_r0_reg_6_inst : dff port map( d => registers_n238, gclk 
                           => clk, rnot => registers_n33, q => 
                           mem_sipo_r0_6_port);
   registers_mem_sipo_r0_reg_7_inst : dff port map( d => registers_n239, gclk 
                           => clk, rnot => registers_n34, q => 
                           mem_sipo_r0_7_port);
   registers_s_mem_sipo_g0_reg_0_inst : dff port map( d => registers_n240, gclk
                           => clk, rnot => registers_n35, q => 
                           registers_s_mem_sipo_g0_0_port);
   registers_s_mem_sipo_g0_reg_1_inst : dff port map( d => registers_n241, gclk
                           => clk, rnot => registers_n36, q => 
                           registers_s_mem_sipo_g0_1_port);
   registers_s_mem_sipo_g0_reg_2_inst : dff port map( d => registers_n242, gclk
                           => clk, rnot => registers_n37, q => 
                           registers_s_mem_sipo_g0_2_port);
   registers_s_mem_sipo_g0_reg_3_inst : dff port map( d => registers_n243, gclk
                           => clk, rnot => registers_n38, q => 
                           registers_s_mem_sipo_g0_3_port);
   registers_s_mem_sipo_g0_reg_4_inst : dff port map( d => registers_n244, gclk
                           => clk, rnot => registers_n39, q => 
                           registers_s_mem_sipo_g0_4_port);
   registers_s_mem_sipo_g0_reg_5_inst : dff port map( d => registers_n245, gclk
                           => clk, rnot => registers_n40, q => 
                           registers_s_mem_sipo_g0_5_port);
   registers_s_mem_sipo_g0_reg_6_inst : dff port map( d => registers_n246, gclk
                           => clk, rnot => registers_n41, q => 
                           registers_s_mem_sipo_g0_6_port);
   registers_s_mem_sipo_g0_reg_7_inst : dff port map( d => registers_n247, gclk
                           => clk, rnot => registers_n42, q => 
                           registers_s_mem_sipo_g0_7_port);
   registers_s_mem_sipo_r0_reg_0_inst : dff port map( d => registers_n248, gclk
                           => clk, rnot => registers_n43, q => 
                           registers_s_mem_sipo_r0_0_port);
   registers_s_mem_sipo_r0_reg_1_inst : dff port map( d => registers_n249, gclk
                           => clk, rnot => registers_n44, q => 
                           registers_s_mem_sipo_r0_1_port);
   registers_s_mem_sipo_r0_reg_2_inst : dff port map( d => registers_n250, gclk
                           => clk, rnot => registers_n45, q => 
                           registers_s_mem_sipo_r0_2_port);
   registers_s_mem_sipo_r0_reg_3_inst : dff port map( d => registers_n251, gclk
                           => clk, rnot => registers_n46, q => 
                           registers_s_mem_sipo_r0_3_port);
   registers_s_mem_sipo_r0_reg_4_inst : dff port map( d => registers_n252, gclk
                           => clk, rnot => registers_n47, q => 
                           registers_s_mem_sipo_r0_4_port);
   registers_s_mem_sipo_r0_reg_5_inst : dff port map( d => registers_n253, gclk
                           => clk, rnot => registers_n48, q => 
                           registers_s_mem_sipo_r0_5_port);
   registers_s_mem_sipo_r0_reg_6_inst : dff port map( d => registers_n254, gclk
                           => clk, rnot => registers_n49, q => 
                           registers_s_mem_sipo_r0_6_port);
   registers_s_mem_sipo_r0_reg_7_inst : dff port map( d => registers_n255, gclk
                           => clk, rnot => registers_n50, q => 
                           registers_s_mem_sipo_r0_7_port);
   registers_mem_sipo_b0_reg_0_inst : dff port map( d => registers_n256, gclk 
                           => clk, rnot => registers_n51, q => 
                           mem_sipo_b0_0_port);
   registers_s_mem_sipo_b0_reg_0_inst : dff port map( d => registers_n257, gclk
                           => clk, rnot => registers_n52, q => 
                           registers_s_mem_sipo_b0_0_port);
   registers_mem_sipo_b0_reg_1_inst : dff port map( d => registers_n258, gclk 
                           => clk, rnot => registers_n53, q => 
                           mem_sipo_b0_1_port);
   registers_s_mem_sipo_b0_reg_1_inst : dff port map( d => registers_n259, gclk
                           => clk, rnot => registers_n54, q => 
                           registers_s_mem_sipo_b0_1_port);
   registers_mem_sipo_b0_reg_2_inst : dff port map( d => registers_n260, gclk 
                           => clk, rnot => registers_n55, q => 
                           mem_sipo_b0_2_port);
   registers_s_mem_sipo_b0_reg_2_inst : dff port map( d => registers_n261, gclk
                           => clk, rnot => registers_n56, q => 
                           registers_s_mem_sipo_b0_2_port);
   registers_mem_sipo_b0_reg_3_inst : dff port map( d => registers_n262, gclk 
                           => clk, rnot => registers_n57, q => 
                           mem_sipo_b0_3_port);
   registers_s_mem_sipo_b0_reg_3_inst : dff port map( d => registers_n263, gclk
                           => clk, rnot => registers_n58, q => 
                           registers_s_mem_sipo_b0_3_port);
   registers_mem_sipo_b0_reg_4_inst : dff port map( d => registers_n264, gclk 
                           => clk, rnot => registers_n59, q => 
                           mem_sipo_b0_4_port);
   registers_s_mem_sipo_b0_reg_4_inst : dff port map( d => registers_n265, gclk
                           => clk, rnot => registers_n60, q => 
                           registers_s_mem_sipo_b0_4_port);
   registers_mem_sipo_b0_reg_5_inst : dff port map( d => registers_n266, gclk 
                           => clk, rnot => registers_n61, q => 
                           mem_sipo_b0_5_port);
   registers_s_mem_sipo_b0_reg_5_inst : dff port map( d => registers_n267, gclk
                           => clk, rnot => registers_n62, q => 
                           registers_s_mem_sipo_b0_5_port);
   registers_mem_sipo_b0_reg_6_inst : dff port map( d => registers_n268, gclk 
                           => clk, rnot => registers_n63, q => 
                           mem_sipo_b0_6_port);
   registers_s_mem_sipo_b0_reg_6_inst : dff port map( d => registers_n269, gclk
                           => clk, rnot => registers_n64, q => 
                           registers_s_mem_sipo_b0_6_port);
   registers_mem_sipo_b0_reg_7_inst : dff port map( d => registers_n270, gclk 
                           => clk, rnot => registers_n65, q => 
                           mem_sipo_b0_7_port);
   registers_s_mem_sipo_b0_reg_7_inst : dff port map( d => registers_n271, gclk
                           => clk, rnot => registers_n66, q => 
                           registers_s_mem_sipo_b0_7_port);
   registers_reg_hub_f_reg : dff port map( d => registers_n272, gclk => clk, 
                           rnot => registers_n67, q => reg_hub_f);
   registers_addr_i_reg_1_inst : dff port map( d => registers_n282, gclk => clk
                           , rnot => registers_n68, q => addr_i_1_port);
   registers_addr_i_reg_2_inst : dff port map( d => registers_n273, gclk => clk
                           , rnot => registers_n69, q => addr_i_2_port);
   registers_addr_i_reg_3_inst : dff port map( d => registers_n275, gclk => clk
                           , rnot => registers_n70, q => addr_i_3_port);
   registers_addr_i_reg_0_inst : dff port map( d => registers_n280, gclk => clk
                           , rnot => registers_n71, q => addr_i_0_port);
   registers_reg_row_reg_1_inst : dff port map( d => registers_n276, gclk => 
                           clk, rnot => registers_n72, q => 
                           registers_reg_row_1_port);
   registers_reg_cd_reg_0_inst : dff port map( d => registers_n278, gclk => clk
                           , rnot => registers_n73, q => 
                           registers_reg_cd_0_port);
   registers_reg_cd_reg_2_inst : dff port map( d => registers_n279, gclk => clk
                           , rnot => registers_n74, q => 
                           registers_reg_cd_2_port);
   registers_reg_cd_reg_1_inst : dff port map( d => registers_n277, gclk => clk
                           , rnot => registers_n75, q => 
                           registers_reg_cd_1_port);
   registers_reg_row_reg_0_inst : dff port map( d => registers_n274, gclk => 
                           clk, rnot => registers_n76, q => 
                           registers_reg_row_0_port);
   registers_mem_to_reg_reg_1_inst : dff port map( d => registers_n284, gclk =>
                           clk, rnot => registers_n77, q => 
                           registers_mem_to_reg_1_port);
   registers_reg_col_inc_reg_0_inst : dff port map( d => registers_n281, gclk 
                           => clk, rnot => registers_n78, q => 
                           registers_reg_col_inc_0_port);
   registers_reg_col_inc_reg_1_inst : dff port map( d => registers_n283, gclk 
                           => clk, rnot => registers_n79, q => 
                           registers_reg_col_inc_1_port);
   registers_mem_to_reg_reg_0_inst : dff port map( d => n1978, gclk => clk, 
                           rnot => registers_n80, q => 
                           registers_mem_to_reg_0_port);
   registers_s_delay_reg_1_inst : dff port map( d => registers_n285, gclk => 
                           clk, rnot => registers_n81, q => 
                           registers_s_delay_1_port);
   registers_s_delay_reg_0_inst : dff port map( d => registers_n286, gclk => 
                           clk, rnot => registers_n82, q => 
                           registers_s_delay_0_port);
   load_n_store_n92 <= '1';
   load_n_store_n91 <= '1';
   load_n_store_n90 <= '1';
   load_n_store_n89 <= '1';
   load_n_store_n88 <= '1';
   load_n_store_n87 <= '1';
   load_n_store_n86 <= '1';
   load_n_store_n85 <= '1';
   load_n_store_n84 <= '1';
   load_n_store_n83 <= '1';
   load_n_store_n82 <= '1';
   load_n_store_n81 <= '1';
   load_n_store_n80 <= '1';
   load_n_store_n79 <= '1';
   load_n_store_n78 <= '1';
   load_n_store_n77 <= '1';
   load_n_store_n76 <= '1';
   load_n_store_n75 <= '1';
   load_n_store_n74 <= '1';
   load_n_store_n73 <= '1';
   load_n_store_n72 <= '1';
   load_n_store_n71 <= '1';
   load_n_store_n70 <= '1';
   load_n_store_n69 <= '1';
   load_n_store_n68 <= '1';
   load_n_store_n67 <= '1';
   load_n_store_n66 <= '1';
   load_n_store_n65 <= '1';
   load_n_store_n64 <= '1';
   load_n_store_n63 <= '1';
   load_n_store_n62 <= '1';
   load_n_store_n61 <= '1';
   load_n_store_n60 <= '1';
   load_n_store_n59 <= '1';
   load_n_store_n58 <= '1';
   load_n_store_n57 <= '1';
   load_n_store_n56 <= '1';
   load_n_store_n55 <= '1';
   load_n_store_n54 <= '1';
   load_n_store_n53 <= '1';
   load_n_store_n52 <= '1';
   load_n_store_n51 <= '1';
   load_n_store_n50 <= '1';
   load_n_store_n49 <= '1';
   load_n_store_n48 <= '1';
   load_n_store_n47 <= '1';
   load_n_store_n46 <= '1';
   load_n_store_n45 <= '1';
   load_n_store_n44 <= '1';
   load_n_store_n43 <= '1';
   load_n_store_n42 <= '1';
   load_n_store_n41 <= '1';
   load_n_store_n40 <= '1';
   load_n_store_n39 <= '1';
   load_n_store_n38 <= '1';
   load_n_store_n37 <= '1';
   load_n_store_n36 <= '1';
   load_n_store_n35 <= '1';
   load_n_store_n34 <= '1';
   load_n_store_n33 <= '1';
   load_n_store_n32 <= '1';
   load_n_store_n31 <= '1';
   load_n_store_n30 <= '1';
   load_n_store_n29 <= '1';
   load_n_store_n28 <= '1';
   load_n_store_n27 <= '1';
   load_n_store_n26 <= '1';
   load_n_store_n25 <= '1';
   load_n_store_n24 <= '1';
   load_n_store_n23 <= '1';
   load_n_store_n22 <= '1';
   load_n_store_n21 <= '1';
   load_n_store_n20 <= '1';
   load_n_store_n19 <= '1';
   load_n_store_n18 <= '1';
   load_n_store_n17 <= '1';
   load_n_store_n16 <= '1';
   load_n_store_n15 <= '1';
   load_n_store_n14 <= '1';
   load_n_store_n13 <= '1';
   load_n_store_n12 <= '1';
   load_n_store_n11 <= '1';
   load_n_store_n10 <= '1';
   load_n_store_n9 <= '1';
   load_n_store_n8 <= '1';
   load_n_store_n7 <= '1';
   load_n_store_mem_out_b0_reg_7_inst : dff port map( d => n1974, gclk => clk, 
                           rnot => load_n_store_n7, q => mem_out_b0_7_port);
   load_n_store_mem_out_b0_reg_6_inst : dff port map( d => n1973, gclk => clk, 
                           rnot => load_n_store_n8, q => mem_out_b0_6_port);
   load_n_store_mem_out_b0_reg_5_inst : dff port map( d => n1972, gclk => clk, 
                           rnot => load_n_store_n9, q => mem_out_b0_5_port);
   load_n_store_mem_out_b0_reg_4_inst : dff port map( d => n1971, gclk => clk, 
                           rnot => load_n_store_n10, q => mem_out_b0_4_port);
   load_n_store_mem_out_b0_reg_3_inst : dff port map( d => n1970, gclk => clk, 
                           rnot => load_n_store_n11, q => mem_out_b0_3_port);
   load_n_store_mem_out_b0_reg_2_inst : dff port map( d => n1969, gclk => clk, 
                           rnot => load_n_store_n12, q => mem_out_b0_2_port);
   load_n_store_mem_out_b0_reg_1_inst : dff port map( d => n1968, gclk => clk, 
                           rnot => load_n_store_n13, q => mem_out_b0_1_port);
   load_n_store_mem_out_b0_reg_0_inst : dff port map( d => n1967, gclk => clk, 
                           rnot => load_n_store_n14, q => mem_out_b0_0_port);
   load_n_store_lazy_in_reg_0_7_inst : dff port map( d => n1918, gclk => clk, 
                           rnot => load_n_store_n15, q => 
                           load_n_store_lazy_in_0_7_port);
   load_n_store_lazy_in_reg_0_6_inst : dff port map( d => n1917, gclk => clk, 
                           rnot => load_n_store_n16, q => 
                           load_n_store_lazy_in_0_6_port);
   load_n_store_lazy_in_reg_0_5_inst : dff port map( d => n1916, gclk => clk, 
                           rnot => load_n_store_n17, q => 
                           load_n_store_lazy_in_0_5_port);
   load_n_store_lazy_in_reg_0_4_inst : dff port map( d => n1915, gclk => clk, 
                           rnot => load_n_store_n18, q => 
                           load_n_store_lazy_in_0_4_port);
   load_n_store_lazy_in_reg_0_3_inst : dff port map( d => n1914, gclk => clk, 
                           rnot => load_n_store_n19, q => 
                           load_n_store_lazy_in_0_3_port);
   load_n_store_lazy_in_reg_0_2_inst : dff port map( d => n1913, gclk => clk, 
                           rnot => load_n_store_n20, q => 
                           load_n_store_lazy_in_0_2_port);
   load_n_store_lazy_in_reg_0_1_inst : dff port map( d => n1912, gclk => clk, 
                           rnot => load_n_store_n21, q => 
                           load_n_store_lazy_in_0_1_port);
   load_n_store_lazy_in_reg_0_0_inst : dff port map( d => n1911, gclk => clk, 
                           rnot => load_n_store_n22, q => 
                           load_n_store_lazy_in_0_0_port);
   load_n_store_mem_out_g0_reg_7_inst : dff port map( d => n1966, gclk => clk, 
                           rnot => load_n_store_n23, q => mem_out_g0_7_port);
   load_n_store_mem_out_g0_reg_6_inst : dff port map( d => n1965, gclk => clk, 
                           rnot => load_n_store_n24, q => mem_out_g0_6_port);
   load_n_store_mem_out_g0_reg_5_inst : dff port map( d => n1964, gclk => clk, 
                           rnot => load_n_store_n25, q => mem_out_g0_5_port);
   load_n_store_mem_out_g0_reg_4_inst : dff port map( d => n1963, gclk => clk, 
                           rnot => load_n_store_n26, q => mem_out_g0_4_port);
   load_n_store_mem_out_g0_reg_3_inst : dff port map( d => n1962, gclk => clk, 
                           rnot => load_n_store_n27, q => mem_out_g0_3_port);
   load_n_store_mem_out_g0_reg_2_inst : dff port map( d => n1961, gclk => clk, 
                           rnot => load_n_store_n28, q => mem_out_g0_2_port);
   load_n_store_mem_out_g0_reg_1_inst : dff port map( d => n1960, gclk => clk, 
                           rnot => load_n_store_n29, q => mem_out_g0_1_port);
   load_n_store_mem_out_g0_reg_0_inst : dff port map( d => n1959, gclk => clk, 
                           rnot => load_n_store_n30, q => mem_out_g0_0_port);
   load_n_store_lazy_in_reg_1_7_inst : dff port map( d => n1910, gclk => clk, 
                           rnot => load_n_store_n31, q => 
                           load_n_store_lazy_in_1_7_port);
   load_n_store_lazy_in_reg_1_6_inst : dff port map( d => n1909, gclk => clk, 
                           rnot => load_n_store_n32, q => 
                           load_n_store_lazy_in_1_6_port);
   load_n_store_lazy_in_reg_1_5_inst : dff port map( d => n1908, gclk => clk, 
                           rnot => load_n_store_n33, q => 
                           load_n_store_lazy_in_1_5_port);
   load_n_store_lazy_in_reg_1_4_inst : dff port map( d => n1907, gclk => clk, 
                           rnot => load_n_store_n34, q => 
                           load_n_store_lazy_in_1_4_port);
   load_n_store_lazy_in_reg_1_3_inst : dff port map( d => n1906, gclk => clk, 
                           rnot => load_n_store_n35, q => 
                           load_n_store_lazy_in_1_3_port);
   load_n_store_lazy_in_reg_1_2_inst : dff port map( d => n1905, gclk => clk, 
                           rnot => load_n_store_n36, q => 
                           load_n_store_lazy_in_1_2_port);
   load_n_store_lazy_in_reg_1_1_inst : dff port map( d => n1904, gclk => clk, 
                           rnot => load_n_store_n37, q => 
                           load_n_store_lazy_in_1_1_port);
   load_n_store_lazy_in_reg_1_0_inst : dff port map( d => n1903, gclk => clk, 
                           rnot => load_n_store_n38, q => 
                           load_n_store_lazy_in_1_0_port);
   load_n_store_mem_out_r0_reg_7_inst : dff port map( d => n1958, gclk => clk, 
                           rnot => load_n_store_n39, q => mem_out_r0_7_port);
   load_n_store_mem_out_r0_reg_6_inst : dff port map( d => n1957, gclk => clk, 
                           rnot => load_n_store_n40, q => mem_out_r0_6_port);
   load_n_store_mem_out_r0_reg_5_inst : dff port map( d => n1956, gclk => clk, 
                           rnot => load_n_store_n41, q => mem_out_r0_5_port);
   load_n_store_mem_out_r0_reg_4_inst : dff port map( d => n1955, gclk => clk, 
                           rnot => load_n_store_n42, q => mem_out_r0_4_port);
   load_n_store_mem_out_r0_reg_3_inst : dff port map( d => n1954, gclk => clk, 
                           rnot => load_n_store_n43, q => mem_out_r0_3_port);
   load_n_store_mem_out_r0_reg_2_inst : dff port map( d => n1953, gclk => clk, 
                           rnot => load_n_store_n44, q => mem_out_r0_2_port);
   load_n_store_mem_out_r0_reg_1_inst : dff port map( d => n1952, gclk => clk, 
                           rnot => load_n_store_n45, q => mem_out_r0_1_port);
   load_n_store_mem_out_r0_reg_0_inst : dff port map( d => n1951, gclk => clk, 
                           rnot => load_n_store_n46, q => mem_out_r0_0_port);
   load_n_store_lazy_in_reg_2_7_inst : dff port map( d => n1902, gclk => clk, 
                           rnot => load_n_store_n47, q => 
                           load_n_store_lazy_in_2_7_port);
   load_n_store_lazy_in_reg_2_6_inst : dff port map( d => n1901, gclk => clk, 
                           rnot => load_n_store_n48, q => 
                           load_n_store_lazy_in_2_6_port);
   load_n_store_lazy_in_reg_2_5_inst : dff port map( d => n1900, gclk => clk, 
                           rnot => load_n_store_n49, q => 
                           load_n_store_lazy_in_2_5_port);
   load_n_store_lazy_in_reg_2_4_inst : dff port map( d => n1899, gclk => clk, 
                           rnot => load_n_store_n50, q => 
                           load_n_store_lazy_in_2_4_port);
   load_n_store_lazy_in_reg_2_3_inst : dff port map( d => n1898, gclk => clk, 
                           rnot => load_n_store_n51, q => 
                           load_n_store_lazy_in_2_3_port);
   load_n_store_lazy_in_reg_2_2_inst : dff port map( d => n1897, gclk => clk, 
                           rnot => load_n_store_n52, q => 
                           load_n_store_lazy_in_2_2_port);
   load_n_store_lazy_in_reg_2_1_inst : dff port map( d => n1896, gclk => clk, 
                           rnot => load_n_store_n53, q => 
                           load_n_store_lazy_in_2_1_port);
   load_n_store_lazy_in_reg_2_0_inst : dff port map( d => n1895, gclk => clk, 
                           rnot => load_n_store_n54, q => 
                           load_n_store_lazy_in_2_0_port);
   load_n_store_top_ack_reg : dff port map( d => load_n_store_n301, gclk => clk
                           , rnot => load_n_store_n55, q => top_ack_port);
   load_n_store_we_i_reg : dff port map( d => n1894, gclk => clk, rnot => 
                           load_n_store_n56, q => load_n_store_we_i);
   load_n_store_mem_hub_f_reg : dff port map( d => load_n_store_n300, gclk => 
                           clk, rnot => load_n_store_n57, q => mem_hub_f);
   load_n_store_mem_reg_f_reg : dff port map( d => load_n_store_n299, gclk => 
                           clk, rnot => load_n_store_n58, q => mem_reg_f);
   load_n_store_simple_mem_sm_reg_1_inst : dff port map( d => load_n_store_n303
                           , gclk => clk, rnot => load_n_store_n59, q => 
                           load_n_store_simple_mem_sm_1_port);
   load_n_store_simple_mem_sm_reg_0_inst : dff port map( d => load_n_store_n302
                           , gclk => clk, rnot => load_n_store_n60, q => 
                           load_n_store_simple_mem_sm_0_port);
   load_n_store_mem_timer_reg_30_inst : dff port map( d => n1950, gclk => clk, 
                           rnot => load_n_store_n61, q => 
                           load_n_store_mem_timer_30_port);
   load_n_store_mem_timer_reg_29_inst : dff port map( d => n1949, gclk => clk, 
                           rnot => load_n_store_n62, q => 
                           load_n_store_mem_timer_29_port);
   load_n_store_mem_timer_reg_28_inst : dff port map( d => n1948, gclk => clk, 
                           rnot => load_n_store_n63, q => 
                           load_n_store_mem_timer_28_port);
   load_n_store_mem_timer_reg_27_inst : dff port map( d => n1947, gclk => clk, 
                           rnot => load_n_store_n64, q => 
                           load_n_store_mem_timer_27_port);
   load_n_store_mem_timer_reg_26_inst : dff port map( d => n1946, gclk => clk, 
                           rnot => load_n_store_n65, q => 
                           load_n_store_mem_timer_26_port);
   load_n_store_mem_timer_reg_25_inst : dff port map( d => n1945, gclk => clk, 
                           rnot => load_n_store_n66, q => 
                           load_n_store_mem_timer_25_port);
   load_n_store_mem_timer_reg_24_inst : dff port map( d => n1944, gclk => clk, 
                           rnot => load_n_store_n67, q => 
                           load_n_store_mem_timer_24_port);
   load_n_store_mem_timer_reg_23_inst : dff port map( d => n1943, gclk => clk, 
                           rnot => load_n_store_n68, q => 
                           load_n_store_mem_timer_23_port);
   load_n_store_mem_timer_reg_22_inst : dff port map( d => n1942, gclk => clk, 
                           rnot => load_n_store_n69, q => 
                           load_n_store_mem_timer_22_port);
   load_n_store_mem_timer_reg_21_inst : dff port map( d => n1941, gclk => clk, 
                           rnot => load_n_store_n70, q => 
                           load_n_store_mem_timer_21_port);
   load_n_store_mem_timer_reg_20_inst : dff port map( d => n1940, gclk => clk, 
                           rnot => load_n_store_n71, q => 
                           load_n_store_mem_timer_20_port);
   load_n_store_mem_timer_reg_19_inst : dff port map( d => n1939, gclk => clk, 
                           rnot => load_n_store_n72, q => 
                           load_n_store_mem_timer_19_port);
   load_n_store_mem_timer_reg_18_inst : dff port map( d => n1938, gclk => clk, 
                           rnot => load_n_store_n73, q => 
                           load_n_store_mem_timer_18_port);
   load_n_store_mem_timer_reg_17_inst : dff port map( d => n1937, gclk => clk, 
                           rnot => load_n_store_n74, q => 
                           load_n_store_mem_timer_17_port);
   load_n_store_mem_timer_reg_16_inst : dff port map( d => n1936, gclk => clk, 
                           rnot => load_n_store_n75, q => 
                           load_n_store_mem_timer_16_port);
   load_n_store_mem_timer_reg_15_inst : dff port map( d => n1935, gclk => clk, 
                           rnot => load_n_store_n76, q => 
                           load_n_store_mem_timer_15_port);
   load_n_store_mem_timer_reg_14_inst : dff port map( d => n1934, gclk => clk, 
                           rnot => load_n_store_n77, q => 
                           load_n_store_mem_timer_14_port);
   load_n_store_mem_timer_reg_13_inst : dff port map( d => n1933, gclk => clk, 
                           rnot => load_n_store_n78, q => 
                           load_n_store_mem_timer_13_port);
   load_n_store_mem_timer_reg_12_inst : dff port map( d => n1932, gclk => clk, 
                           rnot => load_n_store_n79, q => 
                           load_n_store_mem_timer_12_port);
   load_n_store_mem_timer_reg_11_inst : dff port map( d => n1931, gclk => clk, 
                           rnot => load_n_store_n80, q => 
                           load_n_store_mem_timer_11_port);
   load_n_store_mem_timer_reg_10_inst : dff port map( d => n1930, gclk => clk, 
                           rnot => load_n_store_n81, q => 
                           load_n_store_mem_timer_10_port);
   load_n_store_mem_timer_reg_9_inst : dff port map( d => n1929, gclk => clk, 
                           rnot => load_n_store_n82, q => 
                           load_n_store_mem_timer_9_port);
   load_n_store_mem_timer_reg_8_inst : dff port map( d => n1928, gclk => clk, 
                           rnot => load_n_store_n83, q => 
                           load_n_store_mem_timer_8_port);
   load_n_store_mem_timer_reg_7_inst : dff port map( d => n1927, gclk => clk, 
                           rnot => load_n_store_n84, q => 
                           load_n_store_mem_timer_7_port);
   load_n_store_mem_timer_reg_6_inst : dff port map( d => n1926, gclk => clk, 
                           rnot => load_n_store_n85, q => 
                           load_n_store_mem_timer_6_port);
   load_n_store_mem_timer_reg_5_inst : dff port map( d => n1925, gclk => clk, 
                           rnot => load_n_store_n86, q => 
                           load_n_store_mem_timer_5_port);
   load_n_store_mem_timer_reg_4_inst : dff port map( d => n1924, gclk => clk, 
                           rnot => load_n_store_n87, q => 
                           load_n_store_mem_timer_4_port);
   load_n_store_mem_timer_reg_3_inst : dff port map( d => n1923, gclk => clk, 
                           rnot => load_n_store_n88, q => 
                           load_n_store_mem_timer_3_port);
   load_n_store_mem_timer_reg_2_inst : dff port map( d => n1922, gclk => clk, 
                           rnot => load_n_store_n89, q => 
                           load_n_store_mem_timer_2_port);
   load_n_store_mem_timer_reg_1_inst : dff port map( d => n1921, gclk => clk, 
                           rnot => load_n_store_n90, q => 
                           load_n_store_mem_timer_1_port);
   load_n_store_mem_timer_reg_0_inst : dff port map( d => n1920, gclk => clk, 
                           rnot => load_n_store_n91, q => 
                           load_n_store_mem_timer_0_port);
   load_n_store_mem_timer_reg_31_inst : dff port map( d => n1919, gclk => clk, 
                           rnot => load_n_store_n92, q => 
                           load_n_store_mem_timer_31_port);
   display_out_n256 <= '1';
   display_out_n255 <= '1';
   display_out_n254 <= '1';
   display_out_n253 <= '1';
   display_out_n252 <= '1';
   display_out_n251 <= '1';
   display_out_n250 <= '1';
   display_out_n249 <= '1';
   display_out_n248 <= '1';
   display_out_n247 <= '1';
   display_out_n246 <= '1';
   display_out_n245 <= '1';
   display_out_n244 <= '1';
   display_out_n243 <= '1';
   display_out_n242 <= '1';
   display_out_n241 <= '1';
   display_out_n240 <= '1';
   display_out_n239 <= '1';
   display_out_n238 <= '1';
   display_out_n237 <= '1';
   display_out_n236 <= '1';
   display_out_n235 <= '1';
   display_out_n234 <= '1';
   display_out_n233 <= '1';
   display_out_n232 <= '1';
   display_out_n231 <= '1';
   display_out_n230 <= '1';
   display_out_n229 <= '1';
   display_out_n228 <= '1';
   display_out_n227 <= '1';
   display_out_n226 <= '1';
   display_out_n225 <= '1';
   display_out_n224 <= '1';
   display_out_n223 <= '1';
   display_out_n222 <= '1';
   display_out_n221 <= '1';
   display_out_n220 <= '1';
   display_out_n219 <= '1';
   display_out_n218 <= '1';
   display_out_n217 <= '1';
   display_out_n216 <= '1';
   display_out_n215 <= '1';
   display_out_n214 <= '1';
   display_out_n213 <= '1';
   display_out_n212 <= '1';
   display_out_n211 <= '1';
   display_out_n210 <= '1';
   display_out_n209 <= '1';
   display_out_n208 <= '1';
   display_out_n207 <= '1';
   display_out_n206 <= '1';
   display_out_n205 <= '1';
   display_out_n204 <= '1';
   display_out_n203 <= '1';
   display_out_n202 <= '1';
   display_out_n201 <= '1';
   display_out_n200 <= '1';
   display_out_n199 <= '1';
   display_out_n198 <= '1';
   display_out_n197 <= '1';
   display_out_n196 <= '1';
   display_out_n195 <= '1';
   display_out_n194 <= '1';
   display_out_n193 <= '1';
   display_out_n192 <= '1';
   display_out_n191 <= '1';
   display_out_n190 <= '1';
   display_out_n189 <= '1';
   display_out_n188 <= '1';
   display_out_n187 <= '1';
   display_out_n186 <= '1';
   display_out_n185 <= '1';
   display_out_n184 <= '1';
   display_out_n183 <= '1';
   display_out_n182 <= '1';
   display_out_n181 <= '1';
   display_out_n180 <= '1';
   display_out_n179 <= '1';
   display_out_n178 <= '1';
   display_out_n177 <= '1';
   display_out_n176 <= '1';
   display_out_n175 <= '1';
   display_out_n174 <= '1';
   display_out_n173 <= '1';
   display_out_n172 <= '1';
   display_out_n171 <= '1';
   display_out_n170 <= '1';
   display_out_n169 <= '1';
   display_out_n168 <= '1';
   display_out_n167 <= '1';
   display_out_n166 <= '1';
   display_out_n165 <= '1';
   display_out_n164 <= '1';
   display_out_n163 <= '1';
   display_out_n162 <= '1';
   display_out_n161 <= '1';
   display_out_n160 <= '1';
   display_out_n159 <= '1';
   display_out_n158 <= '1';
   display_out_n157 <= '1';
   display_out_n156 <= '1';
   display_out_n155 <= '1';
   display_out_n154 <= '1';
   display_out_n153 <= '1';
   display_out_n152 <= '1';
   display_out_n151 <= '1';
   display_out_n150 <= '1';
   display_out_n149 <= '1';
   display_out_n148 <= '1';
   display_out_n147 <= '1';
   display_out_n146 <= '1';
   display_out_n145 <= '1';
   display_out_n144 <= '1';
   display_out_n143 <= '1';
   display_out_n142 <= '1';
   display_out_n141 <= '1';
   display_out_n140 <= '1';
   display_out_n139 <= '1';
   display_out_n138 <= '1';
   display_out_n137 <= '1';
   display_out_n136 <= '1';
   display_out_n135 <= '1';
   display_out_n134 <= '1';
   display_out_n133 <= '1';
   display_out_n132 <= '1';
   display_out_n131 <= '1';
   display_out_n130 <= '1';
   display_out_n129 <= '1';
   display_out_n128 <= '1';
   display_out_n127 <= '1';
   display_out_n126 <= '1';
   display_out_n125 <= '1';
   display_out_n124 <= '1';
   display_out_n123 <= '1';
   display_out_n122 <= '1';
   display_out_n121 <= '1';
   display_out_n120 <= '1';
   display_out_n119 <= '1';
   display_out_n118 <= '1';
   display_out_n117 <= '1';
   display_out_n116 <= '1';
   display_out_n115 <= '1';
   display_out_n114 <= '1';
   display_out_n113 <= '1';
   display_out_n112 <= '1';
   display_out_n111 <= '1';
   display_out_n110 <= '1';
   display_out_n109 <= '1';
   display_out_n108 <= '1';
   display_out_n107 <= '1';
   display_out_n106 <= '1';
   display_out_n105 <= '1';
   display_out_n104 <= '1';
   display_out_n103 <= '1';
   display_out_n102 <= '1';
   display_out_n101 <= '1';
   display_out_n100 <= '1';
   display_out_n99 <= '1';
   display_out_n98 <= '1';
   display_out_n97 <= '1';
   display_out_n96 <= '1';
   display_out_n95 <= '1';
   display_out_n94 <= '1';
   display_out_n93 <= '1';
   display_out_n92 <= '1';
   display_out_n91 <= '1';
   display_out_n90 <= '1';
   display_out_n89 <= '1';
   display_out_n88 <= '1';
   display_out_hub_b0_o_reg : dff port map( d => display_out_n797, gclk => clk,
                           rnot => display_out_n88, q => hub_b0_o_port);
   display_out_hub_g0_o_reg : dff port map( d => display_out_n798, gclk => clk,
                           rnot => display_out_n89, q => hub_g0_o_port);
   display_out_hub_r0_o_reg : dff port map( d => display_out_n799, gclk => clk,
                           rnot => display_out_n90, q => hub_r0_o_port);
   display_out_hub_piso_b0_reg_0_inst : dff port map( d => display_out_n800, 
                           gclk => clk, rnot => display_out_n91, q => 
                           display_out_hub_piso_b0_0_port);
   display_out_hub_piso_b0_reg_1_inst : dff port map( d => display_out_n806, 
                           gclk => clk, rnot => display_out_n92, q => 
                           display_out_hub_piso_b0_1_port);
   display_out_hub_piso_b0_reg_2_inst : dff port map( d => display_out_n805, 
                           gclk => clk, rnot => display_out_n93, q => 
                           display_out_hub_piso_b0_2_port);
   display_out_hub_piso_b0_reg_3_inst : dff port map( d => display_out_n804, 
                           gclk => clk, rnot => display_out_n94, q => 
                           display_out_hub_piso_b0_3_port);
   display_out_hub_piso_b0_reg_4_inst : dff port map( d => display_out_n803, 
                           gclk => clk, rnot => display_out_n95, q => 
                           display_out_hub_piso_b0_4_port);
   display_out_hub_piso_b0_reg_5_inst : dff port map( d => display_out_n802, 
                           gclk => clk, rnot => display_out_n96, q => 
                           display_out_hub_piso_b0_5_port);
   display_out_hub_piso_b0_reg_6_inst : dff port map( d => display_out_n801, 
                           gclk => clk, rnot => display_out_n97, q => 
                           display_out_hub_piso_b0_6_port);
   display_out_hub_piso_b0_reg_7_inst : dff port map( d => n1977, gclk => clk, 
                           rnot => display_out_n98, q => 
                           display_out_hub_piso_b0_7_port);
   display_out_hub_piso_g0_reg_0_inst : dff port map( d => display_out_n807, 
                           gclk => clk, rnot => display_out_n99, q => 
                           display_out_hub_piso_g0_0_port);
   display_out_hub_piso_g0_reg_1_inst : dff port map( d => display_out_n813, 
                           gclk => clk, rnot => display_out_n100, q => 
                           display_out_hub_piso_g0_1_port);
   display_out_hub_piso_g0_reg_2_inst : dff port map( d => display_out_n812, 
                           gclk => clk, rnot => display_out_n101, q => 
                           display_out_hub_piso_g0_2_port);
   display_out_hub_piso_g0_reg_3_inst : dff port map( d => display_out_n811, 
                           gclk => clk, rnot => display_out_n102, q => 
                           display_out_hub_piso_g0_3_port);
   display_out_hub_piso_g0_reg_4_inst : dff port map( d => display_out_n810, 
                           gclk => clk, rnot => display_out_n103, q => 
                           display_out_hub_piso_g0_4_port);
   display_out_hub_piso_g0_reg_5_inst : dff port map( d => display_out_n809, 
                           gclk => clk, rnot => display_out_n104, q => 
                           display_out_hub_piso_g0_5_port);
   display_out_hub_piso_g0_reg_6_inst : dff port map( d => display_out_n808, 
                           gclk => clk, rnot => display_out_n105, q => 
                           display_out_hub_piso_g0_6_port);
   display_out_hub_piso_g0_reg_7_inst : dff port map( d => n1975, gclk => clk, 
                           rnot => display_out_n106, q => 
                           display_out_hub_piso_g0_7_port);
   display_out_hub_piso_r0_reg_0_inst : dff port map( d => display_out_n814, 
                           gclk => clk, rnot => display_out_n107, q => 
                           display_out_hub_piso_r0_0_port);
   display_out_hub_piso_r0_reg_1_inst : dff port map( d => display_out_n820, 
                           gclk => clk, rnot => display_out_n108, q => 
                           display_out_hub_piso_r0_1_port);
   display_out_hub_piso_r0_reg_2_inst : dff port map( d => display_out_n819, 
                           gclk => clk, rnot => display_out_n109, q => 
                           display_out_hub_piso_r0_2_port);
   display_out_hub_piso_r0_reg_3_inst : dff port map( d => display_out_n818, 
                           gclk => clk, rnot => display_out_n110, q => 
                           display_out_hub_piso_r0_3_port);
   display_out_hub_piso_r0_reg_4_inst : dff port map( d => display_out_n817, 
                           gclk => clk, rnot => display_out_n111, q => 
                           display_out_hub_piso_r0_4_port);
   display_out_hub_piso_r0_reg_5_inst : dff port map( d => display_out_n816, 
                           gclk => clk, rnot => display_out_n112, q => 
                           display_out_hub_piso_r0_5_port);
   display_out_hub_piso_r0_reg_6_inst : dff port map( d => display_out_n815, 
                           gclk => clk, rnot => display_out_n113, q => 
                           display_out_hub_piso_r0_6_port);
   display_out_hub_piso_r0_reg_7_inst : dff port map( d => n1976, gclk => clk, 
                           rnot => display_out_n114, q => 
                           display_out_hub_piso_r0_7_port);
   display_out_hub_reg_f_reg : dff port map( d => display_out_n821, gclk => clk
                           , rnot => display_out_n115, q => hub_reg_f);
   display_out_hub_blank_o_reg : dff port map( d => display_out_n826, gclk => 
                           clk, rnot => display_out_n116, q => hub_blank_o_port
                           );
   display_out_disp_timer_reg_31_inst : dff port map( d => n1979, gclk => clk, 
                           rnot => display_out_n117, q => 
                           display_out_disp_timer_31_port);
   display_out_disp_timer_reg_30_inst : dff port map( d => n2012, gclk => clk, 
                           rnot => display_out_n118, q => 
                           display_out_disp_timer_30_port);
   display_out_disp_timer_reg_29_inst : dff port map( d => n2013, gclk => clk, 
                           rnot => display_out_n119, q => 
                           display_out_disp_timer_29_port);
   display_out_disp_timer_reg_28_inst : dff port map( d => n2014, gclk => clk, 
                           rnot => display_out_n120, q => 
                           display_out_disp_timer_28_port);
   display_out_disp_timer_reg_27_inst : dff port map( d => n2015, gclk => clk, 
                           rnot => display_out_n121, q => 
                           display_out_disp_timer_27_port);
   display_out_disp_timer_reg_26_inst : dff port map( d => n2016, gclk => clk, 
                           rnot => display_out_n122, q => 
                           display_out_disp_timer_26_port);
   display_out_disp_timer_reg_25_inst : dff port map( d => n2017, gclk => clk, 
                           rnot => display_out_n123, q => 
                           display_out_disp_timer_25_port);
   display_out_disp_timer_reg_24_inst : dff port map( d => n2018, gclk => clk, 
                           rnot => display_out_n124, q => 
                           display_out_disp_timer_24_port);
   display_out_disp_timer_reg_23_inst : dff port map( d => n2019, gclk => clk, 
                           rnot => display_out_n125, q => 
                           display_out_disp_timer_23_port);
   display_out_disp_timer_reg_22_inst : dff port map( d => n2020, gclk => clk, 
                           rnot => display_out_n126, q => 
                           display_out_disp_timer_22_port);
   display_out_disp_timer_reg_21_inst : dff port map( d => n2021, gclk => clk, 
                           rnot => display_out_n127, q => 
                           display_out_disp_timer_21_port);
   display_out_disp_timer_reg_20_inst : dff port map( d => n2022, gclk => clk, 
                           rnot => display_out_n128, q => 
                           display_out_disp_timer_20_port);
   display_out_disp_timer_reg_19_inst : dff port map( d => n2023, gclk => clk, 
                           rnot => display_out_n129, q => 
                           display_out_disp_timer_19_port);
   display_out_disp_timer_reg_18_inst : dff port map( d => n2024, gclk => clk, 
                           rnot => display_out_n130, q => 
                           display_out_disp_timer_18_port);
   display_out_disp_timer_reg_17_inst : dff port map( d => n2025, gclk => clk, 
                           rnot => display_out_n131, q => 
                           display_out_disp_timer_17_port);
   display_out_disp_timer_reg_16_inst : dff port map( d => n2026, gclk => clk, 
                           rnot => display_out_n132, q => 
                           display_out_disp_timer_16_port);
   display_out_disp_timer_reg_15_inst : dff port map( d => n2027, gclk => clk, 
                           rnot => display_out_n133, q => 
                           display_out_disp_timer_15_port);
   display_out_disp_timer_reg_14_inst : dff port map( d => n2028, gclk => clk, 
                           rnot => display_out_n134, q => 
                           display_out_disp_timer_14_port);
   display_out_disp_timer_reg_13_inst : dff port map( d => display_out_n839, 
                           gclk => clk, rnot => display_out_n135, q => 
                           display_out_disp_timer_13_port);
   display_out_disp_timer_reg_12_inst : dff port map( d => display_out_n838, 
                           gclk => clk, rnot => display_out_n136, q => 
                           display_out_disp_timer_12_port);
   display_out_disp_timer_reg_11_inst : dff port map( d => display_out_n837, 
                           gclk => clk, rnot => display_out_n137, q => 
                           display_out_disp_timer_11_port);
   display_out_disp_timer_reg_10_inst : dff port map( d => display_out_n836, 
                           gclk => clk, rnot => display_out_n138, q => 
                           display_out_disp_timer_10_port);
   display_out_disp_timer_reg_9_inst : dff port map( d => display_out_n835, 
                           gclk => clk, rnot => display_out_n139, q => 
                           display_out_disp_timer_9_port);
   display_out_disp_timer_reg_8_inst : dff port map( d => display_out_n834, 
                           gclk => clk, rnot => display_out_n140, q => 
                           display_out_disp_timer_8_port);
   display_out_disp_timer_reg_6_inst : dff port map( d => display_out_n832, 
                           gclk => clk, rnot => display_out_n141, q => 
                           display_out_disp_timer_6_port);
   display_out_disp_timer_reg_5_inst : dff port map( d => display_out_n831, 
                           gclk => clk, rnot => display_out_n142, q => 
                           display_out_disp_timer_5_port);
   display_out_disp_timer_reg_4_inst : dff port map( d => display_out_n830, 
                           gclk => clk, rnot => display_out_n143, q => 
                           display_out_disp_timer_4_port);
   display_out_disp_timer_reg_3_inst : dff port map( d => display_out_n829, 
                           gclk => clk, rnot => display_out_n144, q => 
                           display_out_disp_timer_3_port);
   display_out_disp_timer_reg_2_inst : dff port map( d => display_out_n828, 
                           gclk => clk, rnot => display_out_n145, q => 
                           display_out_disp_timer_2_port);
   display_out_disp_timer_reg_0_inst : dff port map( d => display_out_n840, 
                           gclk => clk, rnot => display_out_n146, q => 
                           display_out_disp_timer_0_port);
   display_out_disp_timer_reg_1_inst : dff port map( d => display_out_n827, 
                           gclk => clk, rnot => display_out_n147, q => 
                           display_out_disp_timer_1_port);
   display_out_hub_mux_o_reg_1_inst : dff port map( d => display_out_n824, gclk
                           => clk, rnot => display_out_n148, q => 
                           hub_mux_o_1_port);
   display_out_h_col_reg_31_inst : dff port map( d => display_out_n909, gclk =>
                           clk, rnot => display_out_n149, q => 
                           display_out_h_col_31_port);
   display_out_hub_clk_o_reg : dff port map( d => display_out_n845, gclk => clk
                           , rnot => display_out_n150, q => hub_clk_o_port);
   display_out_clk_timer_reg_2_inst : dff port map( d => display_out_n879, gclk
                           => clk, rnot => display_out_n151, q => 
                           display_out_clk_timer_2_port);
   display_out_clk_timer_reg_3_inst : dff port map( d => display_out_n880, gclk
                           => clk, rnot => display_out_n152, q => 
                           display_out_clk_timer_3_port);
   display_out_clk_timer_reg_4_inst : dff port map( d => display_out_n881, gclk
                           => clk, rnot => display_out_n153, q => 
                           display_out_clk_timer_4_port);
   display_out_clk_timer_reg_0_inst : dff port map( d => display_out_n908, gclk
                           => clk, rnot => display_out_n154, q => 
                           display_out_clk_timer_0_port);
   display_out_clk_timer_reg_30_inst : dff port map( d => display_out_n907, 
                           gclk => clk, rnot => display_out_n155, q => 
                           display_out_clk_timer_30_port);
   display_out_clk_timer_reg_29_inst : dff port map( d => display_out_n906, 
                           gclk => clk, rnot => display_out_n156, q => 
                           display_out_clk_timer_29_port);
   display_out_clk_timer_reg_28_inst : dff port map( d => display_out_n905, 
                           gclk => clk, rnot => display_out_n157, q => 
                           display_out_clk_timer_28_port);
   display_out_clk_timer_reg_27_inst : dff port map( d => display_out_n904, 
                           gclk => clk, rnot => display_out_n158, q => 
                           display_out_clk_timer_27_port);
   display_out_clk_timer_reg_26_inst : dff port map( d => display_out_n903, 
                           gclk => clk, rnot => display_out_n159, q => 
                           display_out_clk_timer_26_port);
   display_out_clk_timer_reg_25_inst : dff port map( d => display_out_n902, 
                           gclk => clk, rnot => display_out_n160, q => 
                           display_out_clk_timer_25_port);
   display_out_clk_timer_reg_24_inst : dff port map( d => display_out_n901, 
                           gclk => clk, rnot => display_out_n161, q => 
                           display_out_clk_timer_24_port);
   display_out_clk_timer_reg_23_inst : dff port map( d => display_out_n900, 
                           gclk => clk, rnot => display_out_n162, q => 
                           display_out_clk_timer_23_port);
   display_out_clk_timer_reg_22_inst : dff port map( d => display_out_n899, 
                           gclk => clk, rnot => display_out_n163, q => 
                           display_out_clk_timer_22_port);
   display_out_clk_timer_reg_21_inst : dff port map( d => display_out_n898, 
                           gclk => clk, rnot => display_out_n164, q => 
                           display_out_clk_timer_21_port);
   display_out_clk_timer_reg_20_inst : dff port map( d => display_out_n897, 
                           gclk => clk, rnot => display_out_n165, q => 
                           display_out_clk_timer_20_port);
   display_out_clk_timer_reg_19_inst : dff port map( d => display_out_n896, 
                           gclk => clk, rnot => display_out_n166, q => 
                           display_out_clk_timer_19_port);
   display_out_clk_timer_reg_18_inst : dff port map( d => display_out_n895, 
                           gclk => clk, rnot => display_out_n167, q => 
                           display_out_clk_timer_18_port);
   display_out_clk_timer_reg_17_inst : dff port map( d => display_out_n894, 
                           gclk => clk, rnot => display_out_n168, q => 
                           display_out_clk_timer_17_port);
   display_out_clk_timer_reg_16_inst : dff port map( d => display_out_n893, 
                           gclk => clk, rnot => display_out_n169, q => 
                           display_out_clk_timer_16_port);
   display_out_clk_timer_reg_15_inst : dff port map( d => display_out_n892, 
                           gclk => clk, rnot => display_out_n170, q => 
                           display_out_clk_timer_15_port);
   display_out_clk_timer_reg_14_inst : dff port map( d => display_out_n891, 
                           gclk => clk, rnot => display_out_n171, q => 
                           display_out_clk_timer_14_port);
   display_out_clk_timer_reg_13_inst : dff port map( d => display_out_n890, 
                           gclk => clk, rnot => display_out_n172, q => 
                           display_out_clk_timer_13_port);
   display_out_clk_timer_reg_12_inst : dff port map( d => display_out_n889, 
                           gclk => clk, rnot => display_out_n173, q => 
                           display_out_clk_timer_12_port);
   display_out_clk_timer_reg_11_inst : dff port map( d => display_out_n888, 
                           gclk => clk, rnot => display_out_n174, q => 
                           display_out_clk_timer_11_port);
   display_out_clk_timer_reg_10_inst : dff port map( d => display_out_n887, 
                           gclk => clk, rnot => display_out_n175, q => 
                           display_out_clk_timer_10_port);
   display_out_clk_timer_reg_9_inst : dff port map( d => display_out_n886, gclk
                           => clk, rnot => display_out_n176, q => 
                           display_out_clk_timer_9_port);
   display_out_clk_timer_reg_8_inst : dff port map( d => display_out_n885, gclk
                           => clk, rnot => display_out_n177, q => 
                           display_out_clk_timer_8_port);
   display_out_clk_timer_reg_7_inst : dff port map( d => display_out_n884, gclk
                           => clk, rnot => display_out_n178, q => 
                           display_out_clk_timer_7_port);
   display_out_clk_timer_reg_6_inst : dff port map( d => display_out_n883, gclk
                           => clk, rnot => display_out_n179, q => 
                           display_out_clk_timer_6_port);
   display_out_clk_timer_reg_5_inst : dff port map( d => display_out_n882, gclk
                           => clk, rnot => display_out_n180, q => 
                           display_out_clk_timer_5_port);
   display_out_clk_timer_reg_1_inst : dff port map( d => display_out_n878, gclk
                           => clk, rnot => display_out_n181, q => 
                           display_out_clk_timer_1_port);
   display_out_h_col_reg_0_inst : dff port map( d => display_out_n876, gclk => 
                           clk, rnot => display_out_n182, q => 
                           display_out_h_col_0_port);
   display_out_h_col_reg_30_inst : dff port map( d => display_out_n875, gclk =>
                           clk, rnot => display_out_n183, q => 
                           display_out_h_col_30_port);
   display_out_h_col_reg_29_inst : dff port map( d => display_out_n874, gclk =>
                           clk, rnot => display_out_n184, q => 
                           display_out_h_col_29_port);
   display_out_h_col_reg_28_inst : dff port map( d => display_out_n873, gclk =>
                           clk, rnot => display_out_n185, q => 
                           display_out_h_col_28_port);
   display_out_h_col_reg_27_inst : dff port map( d => display_out_n872, gclk =>
                           clk, rnot => display_out_n186, q => 
                           display_out_h_col_27_port);
   display_out_h_col_reg_26_inst : dff port map( d => display_out_n871, gclk =>
                           clk, rnot => display_out_n187, q => 
                           display_out_h_col_26_port);
   display_out_h_col_reg_25_inst : dff port map( d => display_out_n870, gclk =>
                           clk, rnot => display_out_n188, q => 
                           display_out_h_col_25_port);
   display_out_h_col_reg_24_inst : dff port map( d => display_out_n869, gclk =>
                           clk, rnot => display_out_n189, q => 
                           display_out_h_col_24_port);
   display_out_h_col_reg_23_inst : dff port map( d => display_out_n868, gclk =>
                           clk, rnot => display_out_n190, q => 
                           display_out_h_col_23_port);
   display_out_h_col_reg_22_inst : dff port map( d => display_out_n867, gclk =>
                           clk, rnot => display_out_n191, q => 
                           display_out_h_col_22_port);
   display_out_h_col_reg_21_inst : dff port map( d => display_out_n866, gclk =>
                           clk, rnot => display_out_n192, q => 
                           display_out_h_col_21_port);
   display_out_h_col_reg_20_inst : dff port map( d => display_out_n865, gclk =>
                           clk, rnot => display_out_n193, q => 
                           display_out_h_col_20_port);
   display_out_h_col_reg_19_inst : dff port map( d => display_out_n864, gclk =>
                           clk, rnot => display_out_n194, q => 
                           display_out_h_col_19_port);
   display_out_h_col_reg_18_inst : dff port map( d => display_out_n863, gclk =>
                           clk, rnot => display_out_n195, q => 
                           display_out_h_col_18_port);
   display_out_h_col_reg_17_inst : dff port map( d => display_out_n862, gclk =>
                           clk, rnot => display_out_n196, q => 
                           display_out_h_col_17_port);
   display_out_h_col_reg_16_inst : dff port map( d => display_out_n861, gclk =>
                           clk, rnot => display_out_n197, q => 
                           display_out_h_col_16_port);
   display_out_h_col_reg_15_inst : dff port map( d => display_out_n860, gclk =>
                           clk, rnot => display_out_n198, q => 
                           display_out_h_col_15_port);
   display_out_h_col_reg_14_inst : dff port map( d => display_out_n859, gclk =>
                           clk, rnot => display_out_n199, q => 
                           display_out_h_col_14_port);
   display_out_h_col_reg_13_inst : dff port map( d => display_out_n858, gclk =>
                           clk, rnot => display_out_n200, q => 
                           display_out_h_col_13_port);
   display_out_h_col_reg_12_inst : dff port map( d => display_out_n857, gclk =>
                           clk, rnot => display_out_n201, q => 
                           display_out_h_col_12_port);
   display_out_h_col_reg_11_inst : dff port map( d => display_out_n856, gclk =>
                           clk, rnot => display_out_n202, q => 
                           display_out_h_col_11_port);
   display_out_h_col_reg_10_inst : dff port map( d => display_out_n855, gclk =>
                           clk, rnot => display_out_n203, q => 
                           display_out_h_col_10_port);
   display_out_h_col_reg_9_inst : dff port map( d => display_out_n854, gclk => 
                           clk, rnot => display_out_n204, q => 
                           display_out_h_col_9_port);
   display_out_h_col_reg_8_inst : dff port map( d => display_out_n853, gclk => 
                           clk, rnot => display_out_n205, q => 
                           display_out_h_col_8_port);
   display_out_h_col_reg_7_inst : dff port map( d => display_out_n852, gclk => 
                           clk, rnot => display_out_n206, q => 
                           display_out_h_col_7_port);
   display_out_h_col_reg_6_inst : dff port map( d => display_out_n851, gclk => 
                           clk, rnot => display_out_n207, q => 
                           display_out_h_col_6_port);
   display_out_h_col_reg_5_inst : dff port map( d => display_out_n850, gclk => 
                           clk, rnot => display_out_n208, q => 
                           display_out_h_col_5_port);
   display_out_h_col_reg_4_inst : dff port map( d => display_out_n849, gclk => 
                           clk, rnot => display_out_n209, q => 
                           display_out_h_col_4_port);
   display_out_h_col_reg_3_inst : dff port map( d => display_out_n848, gclk => 
                           clk, rnot => display_out_n210, q => 
                           display_out_h_col_3_port);
   display_out_h_col_reg_2_inst : dff port map( d => display_out_n847, gclk => 
                           clk, rnot => display_out_n211, q => 
                           display_out_h_col_2_port);
   display_out_h_col_reg_1_inst : dff port map( d => display_out_n846, gclk => 
                           clk, rnot => display_out_n212, q => 
                           display_out_h_col_1_port);
   display_out_clk_timer_reg_31_inst : dff port map( d => display_out_n910, 
                           gclk => clk, rnot => display_out_n213, q => 
                           display_out_clk_timer_31_port);
   display_out_h_row_reg_31_inst : dff port map( d => n2001, gclk => clk, rnot 
                           => display_out_n214, q => display_out_h_row_31_port)
                           ;
   display_out_h_row_reg_30_inst : dff port map( d => n2000, gclk => clk, rnot 
                           => display_out_n215, q => display_out_h_row_30_port)
                           ;
   display_out_h_row_reg_29_inst : dff port map( d => n1999, gclk => clk, rnot 
                           => display_out_n216, q => display_out_h_row_29_port)
                           ;
   display_out_h_row_reg_28_inst : dff port map( d => n1998, gclk => clk, rnot 
                           => display_out_n217, q => display_out_h_row_28_port)
                           ;
   display_out_h_row_reg_27_inst : dff port map( d => n1997, gclk => clk, rnot 
                           => display_out_n218, q => display_out_h_row_27_port)
                           ;
   display_out_h_row_reg_26_inst : dff port map( d => n1996, gclk => clk, rnot 
                           => display_out_n219, q => display_out_h_row_26_port)
                           ;
   display_out_h_row_reg_25_inst : dff port map( d => n1995, gclk => clk, rnot 
                           => display_out_n220, q => display_out_h_row_25_port)
                           ;
   display_out_h_row_reg_24_inst : dff port map( d => n1994, gclk => clk, rnot 
                           => display_out_n221, q => display_out_h_row_24_port)
                           ;
   display_out_h_row_reg_23_inst : dff port map( d => n1993, gclk => clk, rnot 
                           => display_out_n222, q => display_out_h_row_23_port)
                           ;
   display_out_h_row_reg_22_inst : dff port map( d => n1992, gclk => clk, rnot 
                           => display_out_n223, q => display_out_h_row_22_port)
                           ;
   display_out_h_row_reg_21_inst : dff port map( d => n1991, gclk => clk, rnot 
                           => display_out_n224, q => display_out_h_row_21_port)
                           ;
   display_out_h_row_reg_20_inst : dff port map( d => n1990, gclk => clk, rnot 
                           => display_out_n225, q => display_out_h_row_20_port)
                           ;
   display_out_h_row_reg_19_inst : dff port map( d => n1989, gclk => clk, rnot 
                           => display_out_n226, q => display_out_h_row_19_port)
                           ;
   display_out_h_row_reg_18_inst : dff port map( d => n1988, gclk => clk, rnot 
                           => display_out_n227, q => display_out_h_row_18_port)
                           ;
   display_out_h_row_reg_17_inst : dff port map( d => n1987, gclk => clk, rnot 
                           => display_out_n228, q => display_out_h_row_17_port)
                           ;
   display_out_h_row_reg_16_inst : dff port map( d => n1986, gclk => clk, rnot 
                           => display_out_n229, q => display_out_h_row_16_port)
                           ;
   display_out_h_row_reg_15_inst : dff port map( d => n1985, gclk => clk, rnot 
                           => display_out_n230, q => display_out_h_row_15_port)
                           ;
   display_out_h_row_reg_14_inst : dff port map( d => n1984, gclk => clk, rnot 
                           => display_out_n231, q => display_out_h_row_14_port)
                           ;
   display_out_h_row_reg_13_inst : dff port map( d => n1983, gclk => clk, rnot 
                           => display_out_n232, q => display_out_h_row_13_port)
                           ;
   display_out_h_row_reg_12_inst : dff port map( d => n1982, gclk => clk, rnot 
                           => display_out_n233, q => display_out_h_row_12_port)
                           ;
   display_out_h_row_reg_11_inst : dff port map( d => n1981, gclk => clk, rnot 
                           => display_out_n234, q => display_out_h_row_11_port)
                           ;
   display_out_h_row_reg_10_inst : dff port map( d => n1980, gclk => clk, rnot 
                           => display_out_n235, q => display_out_h_row_10_port)
                           ;
   display_out_h_row_reg_9_inst : dff port map( d => n2002, gclk => clk, rnot 
                           => display_out_n236, q => display_out_h_row_9_port);
   display_out_h_row_reg_8_inst : dff port map( d => n2003, gclk => clk, rnot 
                           => display_out_n237, q => display_out_h_row_8_port);
   display_out_h_row_reg_7_inst : dff port map( d => n2004, gclk => clk, rnot 
                           => display_out_n238, q => display_out_h_row_7_port);
   display_out_h_row_reg_6_inst : dff port map( d => n2005, gclk => clk, rnot 
                           => display_out_n239, q => display_out_h_row_6_port);
   display_out_h_row_reg_5_inst : dff port map( d => n2006, gclk => clk, rnot 
                           => display_out_n240, q => display_out_h_row_5_port);
   display_out_h_row_reg_4_inst : dff port map( d => n2007, gclk => clk, rnot 
                           => display_out_n241, q => display_out_h_row_4_port);
   display_out_hub_mux_o_reg_3_inst : dff port map( d => display_out_n822, gclk
                           => clk, rnot => display_out_n242, q => 
                           hub_mux_o_3_port);
   display_out_h_row_reg_3_inst : dff port map( d => n2008, gclk => clk, rnot 
                           => display_out_n243, q => display_out_h_row_3_port);
   display_out_hub_mux_o_reg_2_inst : dff port map( d => display_out_n823, gclk
                           => clk, rnot => display_out_n244, q => 
                           hub_mux_o_2_port);
   display_out_h_row_reg_2_inst : dff port map( d => n2009, gclk => clk, rnot 
                           => display_out_n245, q => display_out_h_row_2_port);
   display_out_hub_mux_o_reg_0_inst : dff port map( d => display_out_n825, gclk
                           => clk, rnot => display_out_n246, q => 
                           hub_mux_o_0_port);
   display_out_h_row_reg_0_inst : dff port map( d => n2010, gclk => clk, rnot 
                           => display_out_n247, q => display_out_h_row_0_port);
   display_out_h_row_reg_1_inst : dff port map( d => n2011, gclk => clk, rnot 
                           => display_out_n248, q => display_out_h_row_1_port);
   display_out_bcd_time_reg_2_inst : dff port map( d => display_out_n841, gclk 
                           => clk, rnot => display_out_n249, q => 
                           display_out_bcd_time_2_port);
   display_out_bcd_time_reg_1_inst : dff port map( d => display_out_n843, gclk 
                           => clk, rnot => display_out_n250, q => 
                           display_out_bcd_time_1_port);
   display_out_bcd_time_reg_0_inst : dff port map( d => display_out_n842, gclk 
                           => clk, rnot => display_out_n251, q => 
                           display_out_bcd_time_0_port);
   display_out_hub_latch_o_reg : dff port map( d => display_out_n844, gclk => 
                           clk, rnot => display_out_n252, q => hub_latch_o_port
                           );
   display_out_disp_timer_reg_7_inst : dff port map( d => display_out_n833, 
                           gclk => clk, rnot => display_out_n253, q => 
                           display_out_disp_timer_7_port);
   display_out_hub_out_sm_reg_2_inst : dff port map( d => display_out_n911, 
                           gclk => clk, rnot => display_out_n254, q => 
                           display_out_hub_out_sm_2_port);
   display_out_hub_out_sm_reg_1_inst : dff port map( d => display_out_n877, 
                           gclk => clk, rnot => display_out_n255, q => 
                           display_out_hub_out_sm_1_port);
   display_out_hub_out_sm_reg_0_inst : dff port map( d => display_out_n912, 
                           gclk => clk, rnot => display_out_n256, q => 
                           display_out_hub_out_sm_0_port);
   load_n_store_RGB_Array_0_n472 <= '1';
   load_n_store_RGB_Array_0_n471 <= '1';
   load_n_store_RGB_Array_0_n470 <= '1';
   load_n_store_RGB_Array_0_n469 <= '1';
   load_n_store_RGB_Array_0_n468 <= '1';
   load_n_store_RGB_Array_0_n467 <= '1';
   load_n_store_RGB_Array_0_n466 <= '1';
   load_n_store_RGB_Array_0_n465 <= '1';
   load_n_store_RGB_Array_0_n464 <= '1';
   load_n_store_RGB_Array_0_n463 <= '1';
   load_n_store_RGB_Array_0_n462 <= '1';
   load_n_store_RGB_Array_0_n461 <= '1';
   load_n_store_RGB_Array_0_n460 <= '1';
   load_n_store_RGB_Array_0_n459 <= '1';
   load_n_store_RGB_Array_0_n458 <= '1';
   load_n_store_RGB_Array_0_n457 <= '1';
   load_n_store_RGB_Array_0_n456 <= '1';
   load_n_store_RGB_Array_0_n455 <= '1';
   load_n_store_RGB_Array_0_n454 <= '1';
   load_n_store_RGB_Array_0_n453 <= '1';
   load_n_store_RGB_Array_0_n452 <= '1';
   load_n_store_RGB_Array_0_n451 <= '1';
   load_n_store_RGB_Array_0_n450 <= '1';
   load_n_store_RGB_Array_0_n449 <= '1';
   load_n_store_RGB_Array_0_n448 <= '1';
   load_n_store_RGB_Array_0_n447 <= '1';
   load_n_store_RGB_Array_0_n446 <= '1';
   load_n_store_RGB_Array_0_n445 <= '1';
   load_n_store_RGB_Array_0_n444 <= '1';
   load_n_store_RGB_Array_0_n443 <= '1';
   load_n_store_RGB_Array_0_n442 <= '1';
   load_n_store_RGB_Array_0_n441 <= '1';
   load_n_store_RGB_Array_0_n440 <= '1';
   load_n_store_RGB_Array_0_n439 <= '1';
   load_n_store_RGB_Array_0_n438 <= '1';
   load_n_store_RGB_Array_0_n437 <= '1';
   load_n_store_RGB_Array_0_n436 <= '1';
   load_n_store_RGB_Array_0_n435 <= '1';
   load_n_store_RGB_Array_0_n434 <= '1';
   load_n_store_RGB_Array_0_n433 <= '1';
   load_n_store_RGB_Array_0_n432 <= '1';
   load_n_store_RGB_Array_0_n431 <= '1';
   load_n_store_RGB_Array_0_n430 <= '1';
   load_n_store_RGB_Array_0_n429 <= '1';
   load_n_store_RGB_Array_0_n428 <= '1';
   load_n_store_RGB_Array_0_n427 <= '1';
   load_n_store_RGB_Array_0_n426 <= '1';
   load_n_store_RGB_Array_0_n425 <= '1';
   load_n_store_RGB_Array_0_n424 <= '1';
   load_n_store_RGB_Array_0_n423 <= '1';
   load_n_store_RGB_Array_0_n422 <= '1';
   load_n_store_RGB_Array_0_n421 <= '1';
   load_n_store_RGB_Array_0_n420 <= '1';
   load_n_store_RGB_Array_0_n419 <= '1';
   load_n_store_RGB_Array_0_n418 <= '1';
   load_n_store_RGB_Array_0_n417 <= '1';
   load_n_store_RGB_Array_0_n416 <= '1';
   load_n_store_RGB_Array_0_n415 <= '1';
   load_n_store_RGB_Array_0_n414 <= '1';
   load_n_store_RGB_Array_0_n413 <= '1';
   load_n_store_RGB_Array_0_n412 <= '1';
   load_n_store_RGB_Array_0_n411 <= '1';
   load_n_store_RGB_Array_0_n410 <= '1';
   load_n_store_RGB_Array_0_n409 <= '1';
   load_n_store_RGB_Array_0_n408 <= '1';
   load_n_store_RGB_Array_0_n407 <= '1';
   load_n_store_RGB_Array_0_n406 <= '1';
   load_n_store_RGB_Array_0_n405 <= '1';
   load_n_store_RGB_Array_0_n404 <= '1';
   load_n_store_RGB_Array_0_n403 <= '1';
   load_n_store_RGB_Array_0_n402 <= '1';
   load_n_store_RGB_Array_0_n401 <= '1';
   load_n_store_RGB_Array_0_n400 <= '1';
   load_n_store_RGB_Array_0_n399 <= '1';
   load_n_store_RGB_Array_0_n398 <= '1';
   load_n_store_RGB_Array_0_n397 <= '1';
   load_n_store_RGB_Array_0_n396 <= '1';
   load_n_store_RGB_Array_0_n395 <= '1';
   load_n_store_RGB_Array_0_n394 <= '1';
   load_n_store_RGB_Array_0_n393 <= '1';
   load_n_store_RGB_Array_0_n392 <= '1';
   load_n_store_RGB_Array_0_n391 <= '1';
   load_n_store_RGB_Array_0_n390 <= '1';
   load_n_store_RGB_Array_0_n389 <= '1';
   load_n_store_RGB_Array_0_n388 <= '1';
   load_n_store_RGB_Array_0_n387 <= '1';
   load_n_store_RGB_Array_0_n386 <= '1';
   load_n_store_RGB_Array_0_n385 <= '1';
   load_n_store_RGB_Array_0_n384 <= '1';
   load_n_store_RGB_Array_0_n383 <= '1';
   load_n_store_RGB_Array_0_n382 <= '1';
   load_n_store_RGB_Array_0_n381 <= '1';
   load_n_store_RGB_Array_0_n380 <= '1';
   load_n_store_RGB_Array_0_n379 <= '1';
   load_n_store_RGB_Array_0_n378 <= '1';
   load_n_store_RGB_Array_0_n377 <= '1';
   load_n_store_RGB_Array_0_n376 <= '1';
   load_n_store_RGB_Array_0_n375 <= '1';
   load_n_store_RGB_Array_0_n374 <= '1';
   load_n_store_RGB_Array_0_n373 <= '1';
   load_n_store_RGB_Array_0_n372 <= '1';
   load_n_store_RGB_Array_0_n371 <= '1';
   load_n_store_RGB_Array_0_n370 <= '1';
   load_n_store_RGB_Array_0_n369 <= '1';
   load_n_store_RGB_Array_0_n368 <= '1';
   load_n_store_RGB_Array_0_n367 <= '1';
   load_n_store_RGB_Array_0_n366 <= '1';
   load_n_store_RGB_Array_0_n365 <= '1';
   load_n_store_RGB_Array_0_n364 <= '1';
   load_n_store_RGB_Array_0_n363 <= '1';
   load_n_store_RGB_Array_0_n362 <= '1';
   load_n_store_RGB_Array_0_n361 <= '1';
   load_n_store_RGB_Array_0_n360 <= '1';
   load_n_store_RGB_Array_0_n359 <= '1';
   load_n_store_RGB_Array_0_n358 <= '1';
   load_n_store_RGB_Array_0_n357 <= '1';
   load_n_store_RGB_Array_0_n356 <= '1';
   load_n_store_RGB_Array_0_n355 <= '1';
   load_n_store_RGB_Array_0_n354 <= '1';
   load_n_store_RGB_Array_0_n353 <= '1';
   load_n_store_RGB_Array_0_n352 <= '1';
   load_n_store_RGB_Array_0_n350 <= '1';
   load_n_store_RGB_Array_0_n349 <= '1';
   load_n_store_RGB_Array_0_n347 <= '1';
   load_n_store_RGB_Array_0_n346 <= '1';
   load_n_store_RGB_Array_0_n344 <= '1';
   load_n_store_RGB_Array_0_n343 <= '1';
   load_n_store_RGB_Array_0_n341 <= '1';
   load_n_store_RGB_Array_0_n340 <= '1';
   load_n_store_RGB_Array_0_n338 <= '1';
   load_n_store_RGB_Array_0_n337 <= '1';
   load_n_store_RGB_Array_0_n335 <= '1';
   load_n_store_RGB_Array_0_n334 <= '1';
   load_n_store_RGB_Array_0_n332 <= '1';
   load_n_store_RGB_Array_0_n331 <= '1';
   load_n_store_RGB_Array_0_n329 <= '1';
   load_n_store_RGB_Array_0_data_out_o_reg_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n2, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n329, q => 
                           load_n_store_lazy_out_0_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_0_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n473, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n331, q => 
                           load_n_store_RGB_Array_0_block_ram_r_0_0_port);
   load_n_store_RGB_Array_0_data_out_o_reg_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n36, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n332, q => 
                           load_n_store_lazy_out_0_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_0_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n474, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n334, q => 
                           load_n_store_RGB_Array_0_block_ram_r_0_1_port);
   load_n_store_RGB_Array_0_data_out_o_reg_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n59, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n335, q => 
                           load_n_store_lazy_out_0_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_0_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n475, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n337, q => 
                           load_n_store_RGB_Array_0_block_ram_r_0_2_port);
   load_n_store_RGB_Array_0_data_out_o_reg_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n82, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n338, q => 
                           load_n_store_lazy_out_0_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_0_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n476, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n340, q => 
                           load_n_store_RGB_Array_0_block_ram_r_0_3_port);
   load_n_store_RGB_Array_0_data_out_o_reg_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n105, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n341, q => 
                           load_n_store_lazy_out_0_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_0_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n477, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n343, q => 
                           load_n_store_RGB_Array_0_block_ram_r_0_4_port);
   load_n_store_RGB_Array_0_data_out_o_reg_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n128, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n344, q => 
                           load_n_store_lazy_out_0_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_0_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n478, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n346, q => 
                           load_n_store_RGB_Array_0_block_ram_r_0_5_port);
   load_n_store_RGB_Array_0_data_out_o_reg_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n151, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n347, q => 
                           load_n_store_lazy_out_0_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_0_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n479, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n349, q => 
                           load_n_store_RGB_Array_0_block_ram_r_0_6_port);
   load_n_store_RGB_Array_0_data_out_o_reg_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n174, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n350, q => 
                           load_n_store_lazy_out_0_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_0_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n480, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n352, q => 
                           load_n_store_RGB_Array_0_block_ram_r_0_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_1_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n481, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n353, q => 
                           load_n_store_RGB_Array_0_block_ram_r_1_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_1_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n482, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n354, q => 
                           load_n_store_RGB_Array_0_block_ram_r_1_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_1_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n483, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n355, q => 
                           load_n_store_RGB_Array_0_block_ram_r_1_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_1_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n484, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n356, q => 
                           load_n_store_RGB_Array_0_block_ram_r_1_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_1_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n485, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n357, q => 
                           load_n_store_RGB_Array_0_block_ram_r_1_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_1_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n486, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n358, q => 
                           load_n_store_RGB_Array_0_block_ram_r_1_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_1_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n487, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n359, q => 
                           load_n_store_RGB_Array_0_block_ram_r_1_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_1_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n488, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n360, q => 
                           load_n_store_RGB_Array_0_block_ram_r_1_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_2_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n489, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n361, q => 
                           load_n_store_RGB_Array_0_block_ram_r_2_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_2_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n490, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n362, q => 
                           load_n_store_RGB_Array_0_block_ram_r_2_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_2_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n491, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n363, q => 
                           load_n_store_RGB_Array_0_block_ram_r_2_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_2_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n492, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n364, q => 
                           load_n_store_RGB_Array_0_block_ram_r_2_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_2_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n493, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n365, q => 
                           load_n_store_RGB_Array_0_block_ram_r_2_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_2_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n494, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n366, q => 
                           load_n_store_RGB_Array_0_block_ram_r_2_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_2_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n495, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n367, q => 
                           load_n_store_RGB_Array_0_block_ram_r_2_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_2_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n496, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n368, q => 
                           load_n_store_RGB_Array_0_block_ram_r_2_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_3_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n497, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n369, q => 
                           load_n_store_RGB_Array_0_block_ram_r_3_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_3_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n498, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n370, q => 
                           load_n_store_RGB_Array_0_block_ram_r_3_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_3_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n499, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n371, q => 
                           load_n_store_RGB_Array_0_block_ram_r_3_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_3_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n500, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n372, q => 
                           load_n_store_RGB_Array_0_block_ram_r_3_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_3_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n501, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n373, q => 
                           load_n_store_RGB_Array_0_block_ram_r_3_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_3_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n502, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n374, q => 
                           load_n_store_RGB_Array_0_block_ram_r_3_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_3_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n503, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n375, q => 
                           load_n_store_RGB_Array_0_block_ram_r_3_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_3_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n504, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n376, q => 
                           load_n_store_RGB_Array_0_block_ram_r_3_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_4_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n505, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n377, q => 
                           load_n_store_RGB_Array_0_block_ram_r_4_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_4_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n506, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n378, q => 
                           load_n_store_RGB_Array_0_block_ram_r_4_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_4_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n507, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n379, q => 
                           load_n_store_RGB_Array_0_block_ram_r_4_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_4_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n508, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n380, q => 
                           load_n_store_RGB_Array_0_block_ram_r_4_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_4_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n509, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n381, q => 
                           load_n_store_RGB_Array_0_block_ram_r_4_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_4_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n510, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n382, q => 
                           load_n_store_RGB_Array_0_block_ram_r_4_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_4_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n511, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n383, q => 
                           load_n_store_RGB_Array_0_block_ram_r_4_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_4_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n512, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n384, q => 
                           load_n_store_RGB_Array_0_block_ram_r_4_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_5_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n513, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n385, q => 
                           load_n_store_RGB_Array_0_block_ram_r_5_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_5_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n514, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n386, q => 
                           load_n_store_RGB_Array_0_block_ram_r_5_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_5_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n515, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n387, q => 
                           load_n_store_RGB_Array_0_block_ram_r_5_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_5_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n516, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n388, q => 
                           load_n_store_RGB_Array_0_block_ram_r_5_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_5_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n517, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n389, q => 
                           load_n_store_RGB_Array_0_block_ram_r_5_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_5_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n518, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n390, q => 
                           load_n_store_RGB_Array_0_block_ram_r_5_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_5_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n519, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n391, q => 
                           load_n_store_RGB_Array_0_block_ram_r_5_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_5_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n520, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n392, q => 
                           load_n_store_RGB_Array_0_block_ram_r_5_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_6_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n521, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n393, q => 
                           load_n_store_RGB_Array_0_block_ram_r_6_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_6_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n522, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n394, q => 
                           load_n_store_RGB_Array_0_block_ram_r_6_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_6_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n523, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n395, q => 
                           load_n_store_RGB_Array_0_block_ram_r_6_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_6_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n524, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n396, q => 
                           load_n_store_RGB_Array_0_block_ram_r_6_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_6_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n525, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n397, q => 
                           load_n_store_RGB_Array_0_block_ram_r_6_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_6_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n526, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n398, q => 
                           load_n_store_RGB_Array_0_block_ram_r_6_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_6_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n527, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n399, q => 
                           load_n_store_RGB_Array_0_block_ram_r_6_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_6_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n528, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n400, q => 
                           load_n_store_RGB_Array_0_block_ram_r_6_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_7_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n529, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n401, q => 
                           load_n_store_RGB_Array_0_block_ram_r_7_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_7_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n530, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n402, q => 
                           load_n_store_RGB_Array_0_block_ram_r_7_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_7_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n531, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n403, q => 
                           load_n_store_RGB_Array_0_block_ram_r_7_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_7_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n532, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n404, q => 
                           load_n_store_RGB_Array_0_block_ram_r_7_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_7_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n533, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n405, q => 
                           load_n_store_RGB_Array_0_block_ram_r_7_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_7_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n534, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n406, q => 
                           load_n_store_RGB_Array_0_block_ram_r_7_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_7_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n535, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n407, q => 
                           load_n_store_RGB_Array_0_block_ram_r_7_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_7_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n536, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n408, q => 
                           load_n_store_RGB_Array_0_block_ram_r_7_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_8_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n537, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n409, q => 
                           load_n_store_RGB_Array_0_block_ram_r_8_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_8_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n538, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n410, q => 
                           load_n_store_RGB_Array_0_block_ram_r_8_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_8_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n539, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n411, q => 
                           load_n_store_RGB_Array_0_block_ram_r_8_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_8_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n540, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n412, q => 
                           load_n_store_RGB_Array_0_block_ram_r_8_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_8_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n541, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n413, q => 
                           load_n_store_RGB_Array_0_block_ram_r_8_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_8_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n542, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n414, q => 
                           load_n_store_RGB_Array_0_block_ram_r_8_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_8_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n543, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n415, q => 
                           load_n_store_RGB_Array_0_block_ram_r_8_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_8_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n544, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n416, q => 
                           load_n_store_RGB_Array_0_block_ram_r_8_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_9_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n545, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n417, q => 
                           load_n_store_RGB_Array_0_block_ram_r_9_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_9_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n546, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n418, q => 
                           load_n_store_RGB_Array_0_block_ram_r_9_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_9_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n547, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n419, q => 
                           load_n_store_RGB_Array_0_block_ram_r_9_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_9_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n548, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n420, q => 
                           load_n_store_RGB_Array_0_block_ram_r_9_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_9_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n549, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n421, q => 
                           load_n_store_RGB_Array_0_block_ram_r_9_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_9_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n550, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n422, q => 
                           load_n_store_RGB_Array_0_block_ram_r_9_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_9_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n551, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n423, q => 
                           load_n_store_RGB_Array_0_block_ram_r_9_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_9_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n552, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n424, q => 
                           load_n_store_RGB_Array_0_block_ram_r_9_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_10_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n553, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n425, q => 
                           load_n_store_RGB_Array_0_block_ram_r_10_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_10_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n554, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n426, q => 
                           load_n_store_RGB_Array_0_block_ram_r_10_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_10_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n555, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n427, q => 
                           load_n_store_RGB_Array_0_block_ram_r_10_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_10_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n556, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n428, q => 
                           load_n_store_RGB_Array_0_block_ram_r_10_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_10_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n557, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n429, q => 
                           load_n_store_RGB_Array_0_block_ram_r_10_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_10_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n558, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n430, q => 
                           load_n_store_RGB_Array_0_block_ram_r_10_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_10_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n559, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n431, q => 
                           load_n_store_RGB_Array_0_block_ram_r_10_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_10_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n560, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n432, q => 
                           load_n_store_RGB_Array_0_block_ram_r_10_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_11_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n561, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n433, q => 
                           load_n_store_RGB_Array_0_block_ram_r_11_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_11_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n562, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n434, q => 
                           load_n_store_RGB_Array_0_block_ram_r_11_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_11_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n563, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n435, q => 
                           load_n_store_RGB_Array_0_block_ram_r_11_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_11_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n564, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n436, q => 
                           load_n_store_RGB_Array_0_block_ram_r_11_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_11_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n565, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n437, q => 
                           load_n_store_RGB_Array_0_block_ram_r_11_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_11_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n566, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n438, q => 
                           load_n_store_RGB_Array_0_block_ram_r_11_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_11_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n567, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n439, q => 
                           load_n_store_RGB_Array_0_block_ram_r_11_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_11_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n568, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n440, q => 
                           load_n_store_RGB_Array_0_block_ram_r_11_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_12_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n569, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n441, q => 
                           load_n_store_RGB_Array_0_block_ram_r_12_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_12_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n570, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n442, q => 
                           load_n_store_RGB_Array_0_block_ram_r_12_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_12_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n571, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n443, q => 
                           load_n_store_RGB_Array_0_block_ram_r_12_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_12_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n572, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n444, q => 
                           load_n_store_RGB_Array_0_block_ram_r_12_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_12_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n573, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n445, q => 
                           load_n_store_RGB_Array_0_block_ram_r_12_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_12_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n574, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n446, q => 
                           load_n_store_RGB_Array_0_block_ram_r_12_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_12_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n575, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n447, q => 
                           load_n_store_RGB_Array_0_block_ram_r_12_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_12_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n576, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n448, q => 
                           load_n_store_RGB_Array_0_block_ram_r_12_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_13_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n577, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n449, q => 
                           load_n_store_RGB_Array_0_block_ram_r_13_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_13_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n578, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n450, q => 
                           load_n_store_RGB_Array_0_block_ram_r_13_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_13_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n579, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n451, q => 
                           load_n_store_RGB_Array_0_block_ram_r_13_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_13_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n580, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n452, q => 
                           load_n_store_RGB_Array_0_block_ram_r_13_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_13_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n581, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n453, q => 
                           load_n_store_RGB_Array_0_block_ram_r_13_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_13_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n582, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n454, q => 
                           load_n_store_RGB_Array_0_block_ram_r_13_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_13_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n583, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n455, q => 
                           load_n_store_RGB_Array_0_block_ram_r_13_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_13_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n584, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n456, q => 
                           load_n_store_RGB_Array_0_block_ram_r_13_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_14_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n585, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n457, q => 
                           load_n_store_RGB_Array_0_block_ram_r_14_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_14_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n586, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n458, q => 
                           load_n_store_RGB_Array_0_block_ram_r_14_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_14_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n587, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n459, q => 
                           load_n_store_RGB_Array_0_block_ram_r_14_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_14_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n588, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n460, q => 
                           load_n_store_RGB_Array_0_block_ram_r_14_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_14_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n589, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n461, q => 
                           load_n_store_RGB_Array_0_block_ram_r_14_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_14_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n590, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n462, q => 
                           load_n_store_RGB_Array_0_block_ram_r_14_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_14_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n591, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n463, q => 
                           load_n_store_RGB_Array_0_block_ram_r_14_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_14_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n592, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n464, q => 
                           load_n_store_RGB_Array_0_block_ram_r_14_7_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_15_0_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n593, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n465, q => 
                           load_n_store_RGB_Array_0_block_ram_r_15_0_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_15_1_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n594, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n466, q => 
                           load_n_store_RGB_Array_0_block_ram_r_15_1_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_15_2_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n595, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n467, q => 
                           load_n_store_RGB_Array_0_block_ram_r_15_2_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_15_3_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n596, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n468, q => 
                           load_n_store_RGB_Array_0_block_ram_r_15_3_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_15_4_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n597, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n469, q => 
                           load_n_store_RGB_Array_0_block_ram_r_15_4_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_15_5_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n598, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n470, q => 
                           load_n_store_RGB_Array_0_block_ram_r_15_5_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_15_6_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n599, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n471, q => 
                           load_n_store_RGB_Array_0_block_ram_r_15_6_port);
   load_n_store_RGB_Array_0_block_ram_r_reg_15_7_inst : dff port map( d => 
                           load_n_store_RGB_Array_0_n600, gclk => clk, rnot => 
                           load_n_store_RGB_Array_0_n472, q => 
                           load_n_store_RGB_Array_0_block_ram_r_15_7_port);
   n2444 <= '1';
   n2443 <= '1';
   n2442 <= '1';
   n2441 <= '1';
   n2440 <= '1';
   n2439 <= '1';
   n2438 <= '1';
   n2437 <= '1';
   n2436 <= '1';
   n2435 <= '1';
   n2434 <= '1';
   n2433 <= '1';
   n2432 <= '1';
   n2431 <= '1';
   n2430 <= '1';
   n2429 <= '1';
   n2428 <= '1';
   n2427 <= '1';
   n2426 <= '1';
   n2425 <= '1';
   n2424 <= '1';
   n2423 <= '1';
   n2422 <= '1';
   n2421 <= '1';
   n2420 <= '1';
   n2419 <= '1';
   n2418 <= '1';
   n2417 <= '1';
   n2416 <= '1';
   n2415 <= '1';
   n2414 <= '1';
   n2413 <= '1';
   n2412 <= '1';
   n2411 <= '1';
   n2410 <= '1';
   n2409 <= '1';
   n2408 <= '1';
   n2407 <= '1';
   n2406 <= '1';
   n2405 <= '1';
   n2404 <= '1';
   n2403 <= '1';
   n2402 <= '1';
   n2401 <= '1';
   n2400 <= '1';
   n2399 <= '1';
   n2398 <= '1';
   n2397 <= '1';
   n2396 <= '1';
   n2395 <= '1';
   n2394 <= '1';
   n2393 <= '1';
   n2392 <= '1';
   n2391 <= '1';
   n2390 <= '1';
   n2389 <= '1';
   n2388 <= '1';
   n2387 <= '1';
   n2386 <= '1';
   n2385 <= '1';
   n2384 <= '1';
   n2383 <= '1';
   n2382 <= '1';
   n2381 <= '1';
   n2380 <= '1';
   n2379 <= '1';
   n2378 <= '1';
   n2377 <= '1';
   n2376 <= '1';
   n2375 <= '1';
   n2374 <= '1';
   n2373 <= '1';
   n2372 <= '1';
   n2371 <= '1';
   n2370 <= '1';
   n2369 <= '1';
   n2368 <= '1';
   n2367 <= '1';
   n2366 <= '1';
   n2365 <= '1';
   n2364 <= '1';
   n2363 <= '1';
   n2362 <= '1';
   n2361 <= '1';
   n2360 <= '1';
   n2359 <= '1';
   n2358 <= '1';
   n2357 <= '1';
   n2356 <= '1';
   n2355 <= '1';
   n2354 <= '1';
   n2353 <= '1';
   n2352 <= '1';
   n2351 <= '1';
   n2350 <= '1';
   n2349 <= '1';
   n2348 <= '1';
   n2347 <= '1';
   n2346 <= '1';
   n2345 <= '1';
   n2344 <= '1';
   n2343 <= '1';
   n2342 <= '1';
   n2341 <= '1';
   n2340 <= '1';
   n2339 <= '1';
   n2338 <= '1';
   n2337 <= '1';
   n2336 <= '1';
   n2335 <= '1';
   n2334 <= '1';
   n2333 <= '1';
   n2332 <= '1';
   n2331 <= '1';
   n2330 <= '1';
   n2329 <= '1';
   n2328 <= '1';
   n2327 <= '1';
   n2326 <= '1';
   n2325 <= '1';
   n2324 <= '1';
   n2323 <= '1';
   n2322 <= '1';
   n2321 <= '1';
   n2320 <= '1';
   n2319 <= '1';
   n2318 <= '1';
   n2317 <= '1';
   n2316 <= '1';
   n2315 <= '1';
   n2314 <= '1';
   n2313 <= '1';
   n2312 <= '1';
   n2311 <= '1';
   n2310 <= '1';
   n2309 <= '1';
   load_n_store_RGB_Array_2_data_out_o_reg_0_inst : dff port map( d => n2301, 
                           gclk => clk, rnot => n2309, q => 
                           load_n_store_lazy_out_2_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_0_0_inst : dff port map( d => n2445
                           , gclk => clk, rnot => n2310, q => 
                           load_n_store_RGB_Array_2_block_ram_r_0_0_port);
   load_n_store_RGB_Array_2_data_out_o_reg_1_inst : dff port map( d => n2302, 
                           gclk => clk, rnot => n2311, q => 
                           load_n_store_lazy_out_2_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_0_1_inst : dff port map( d => n2446
                           , gclk => clk, rnot => n2312, q => 
                           load_n_store_RGB_Array_2_block_ram_r_0_1_port);
   load_n_store_RGB_Array_2_data_out_o_reg_2_inst : dff port map( d => n2303, 
                           gclk => clk, rnot => n2313, q => 
                           load_n_store_lazy_out_2_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_0_2_inst : dff port map( d => n2447
                           , gclk => clk, rnot => n2314, q => 
                           load_n_store_RGB_Array_2_block_ram_r_0_2_port);
   load_n_store_RGB_Array_2_data_out_o_reg_3_inst : dff port map( d => n2304, 
                           gclk => clk, rnot => n2315, q => 
                           load_n_store_lazy_out_2_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_0_3_inst : dff port map( d => n2448
                           , gclk => clk, rnot => n2316, q => 
                           load_n_store_RGB_Array_2_block_ram_r_0_3_port);
   load_n_store_RGB_Array_2_data_out_o_reg_4_inst : dff port map( d => n2305, 
                           gclk => clk, rnot => n2317, q => 
                           load_n_store_lazy_out_2_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_0_4_inst : dff port map( d => n2449
                           , gclk => clk, rnot => n2318, q => 
                           load_n_store_RGB_Array_2_block_ram_r_0_4_port);
   load_n_store_RGB_Array_2_data_out_o_reg_5_inst : dff port map( d => n2306, 
                           gclk => clk, rnot => n2319, q => 
                           load_n_store_lazy_out_2_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_0_5_inst : dff port map( d => n2450
                           , gclk => clk, rnot => n2320, q => 
                           load_n_store_RGB_Array_2_block_ram_r_0_5_port);
   load_n_store_RGB_Array_2_data_out_o_reg_6_inst : dff port map( d => n2307, 
                           gclk => clk, rnot => n2321, q => 
                           load_n_store_lazy_out_2_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_0_6_inst : dff port map( d => n2451
                           , gclk => clk, rnot => n2322, q => 
                           load_n_store_RGB_Array_2_block_ram_r_0_6_port);
   load_n_store_RGB_Array_2_data_out_o_reg_7_inst : dff port map( d => n2308, 
                           gclk => clk, rnot => n2323, q => 
                           load_n_store_lazy_out_2_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_0_7_inst : dff port map( d => n2452
                           , gclk => clk, rnot => n2324, q => 
                           load_n_store_RGB_Array_2_block_ram_r_0_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_1_0_inst : dff port map( d => n2453
                           , gclk => clk, rnot => n2325, q => 
                           load_n_store_RGB_Array_2_block_ram_r_1_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_1_1_inst : dff port map( d => n2454
                           , gclk => clk, rnot => n2326, q => 
                           load_n_store_RGB_Array_2_block_ram_r_1_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_1_2_inst : dff port map( d => n2455
                           , gclk => clk, rnot => n2327, q => 
                           load_n_store_RGB_Array_2_block_ram_r_1_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_1_3_inst : dff port map( d => n2456
                           , gclk => clk, rnot => n2328, q => 
                           load_n_store_RGB_Array_2_block_ram_r_1_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_1_4_inst : dff port map( d => n2457
                           , gclk => clk, rnot => n2329, q => 
                           load_n_store_RGB_Array_2_block_ram_r_1_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_1_5_inst : dff port map( d => n2458
                           , gclk => clk, rnot => n2330, q => 
                           load_n_store_RGB_Array_2_block_ram_r_1_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_1_6_inst : dff port map( d => n2459
                           , gclk => clk, rnot => n2331, q => 
                           load_n_store_RGB_Array_2_block_ram_r_1_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_1_7_inst : dff port map( d => n2460
                           , gclk => clk, rnot => n2332, q => 
                           load_n_store_RGB_Array_2_block_ram_r_1_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_2_0_inst : dff port map( d => n2461
                           , gclk => clk, rnot => n2333, q => 
                           load_n_store_RGB_Array_2_block_ram_r_2_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_2_1_inst : dff port map( d => n2462
                           , gclk => clk, rnot => n2334, q => 
                           load_n_store_RGB_Array_2_block_ram_r_2_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_2_2_inst : dff port map( d => n2463
                           , gclk => clk, rnot => n2335, q => 
                           load_n_store_RGB_Array_2_block_ram_r_2_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_2_3_inst : dff port map( d => n2464
                           , gclk => clk, rnot => n2336, q => 
                           load_n_store_RGB_Array_2_block_ram_r_2_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_2_4_inst : dff port map( d => n2465
                           , gclk => clk, rnot => n2337, q => 
                           load_n_store_RGB_Array_2_block_ram_r_2_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_2_5_inst : dff port map( d => n2466
                           , gclk => clk, rnot => n2338, q => 
                           load_n_store_RGB_Array_2_block_ram_r_2_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_2_6_inst : dff port map( d => n2467
                           , gclk => clk, rnot => n2339, q => 
                           load_n_store_RGB_Array_2_block_ram_r_2_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_2_7_inst : dff port map( d => n2468
                           , gclk => clk, rnot => n2340, q => 
                           load_n_store_RGB_Array_2_block_ram_r_2_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_3_0_inst : dff port map( d => n2469
                           , gclk => clk, rnot => n2341, q => 
                           load_n_store_RGB_Array_2_block_ram_r_3_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_3_1_inst : dff port map( d => n2470
                           , gclk => clk, rnot => n2342, q => 
                           load_n_store_RGB_Array_2_block_ram_r_3_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_3_2_inst : dff port map( d => n2471
                           , gclk => clk, rnot => n2343, q => 
                           load_n_store_RGB_Array_2_block_ram_r_3_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_3_3_inst : dff port map( d => n2472
                           , gclk => clk, rnot => n2344, q => 
                           load_n_store_RGB_Array_2_block_ram_r_3_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_3_4_inst : dff port map( d => n2473
                           , gclk => clk, rnot => n2345, q => 
                           load_n_store_RGB_Array_2_block_ram_r_3_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_3_5_inst : dff port map( d => n2474
                           , gclk => clk, rnot => n2346, q => 
                           load_n_store_RGB_Array_2_block_ram_r_3_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_3_6_inst : dff port map( d => n2475
                           , gclk => clk, rnot => n2347, q => 
                           load_n_store_RGB_Array_2_block_ram_r_3_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_3_7_inst : dff port map( d => n2476
                           , gclk => clk, rnot => n2348, q => 
                           load_n_store_RGB_Array_2_block_ram_r_3_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_4_0_inst : dff port map( d => n2477
                           , gclk => clk, rnot => n2349, q => 
                           load_n_store_RGB_Array_2_block_ram_r_4_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_4_1_inst : dff port map( d => n2478
                           , gclk => clk, rnot => n2350, q => 
                           load_n_store_RGB_Array_2_block_ram_r_4_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_4_2_inst : dff port map( d => n2479
                           , gclk => clk, rnot => n2351, q => 
                           load_n_store_RGB_Array_2_block_ram_r_4_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_4_3_inst : dff port map( d => n2480
                           , gclk => clk, rnot => n2352, q => 
                           load_n_store_RGB_Array_2_block_ram_r_4_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_4_4_inst : dff port map( d => n2481
                           , gclk => clk, rnot => n2353, q => 
                           load_n_store_RGB_Array_2_block_ram_r_4_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_4_5_inst : dff port map( d => n2482
                           , gclk => clk, rnot => n2354, q => 
                           load_n_store_RGB_Array_2_block_ram_r_4_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_4_6_inst : dff port map( d => n2483
                           , gclk => clk, rnot => n2355, q => 
                           load_n_store_RGB_Array_2_block_ram_r_4_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_4_7_inst : dff port map( d => n2484
                           , gclk => clk, rnot => n2356, q => 
                           load_n_store_RGB_Array_2_block_ram_r_4_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_5_0_inst : dff port map( d => n2485
                           , gclk => clk, rnot => n2357, q => 
                           load_n_store_RGB_Array_2_block_ram_r_5_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_5_1_inst : dff port map( d => n2486
                           , gclk => clk, rnot => n2358, q => 
                           load_n_store_RGB_Array_2_block_ram_r_5_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_5_2_inst : dff port map( d => n2487
                           , gclk => clk, rnot => n2359, q => 
                           load_n_store_RGB_Array_2_block_ram_r_5_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_5_3_inst : dff port map( d => n2488
                           , gclk => clk, rnot => n2360, q => 
                           load_n_store_RGB_Array_2_block_ram_r_5_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_5_4_inst : dff port map( d => n2489
                           , gclk => clk, rnot => n2361, q => 
                           load_n_store_RGB_Array_2_block_ram_r_5_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_5_5_inst : dff port map( d => n2490
                           , gclk => clk, rnot => n2362, q => 
                           load_n_store_RGB_Array_2_block_ram_r_5_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_5_6_inst : dff port map( d => n2491
                           , gclk => clk, rnot => n2363, q => 
                           load_n_store_RGB_Array_2_block_ram_r_5_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_5_7_inst : dff port map( d => n2492
                           , gclk => clk, rnot => n2364, q => 
                           load_n_store_RGB_Array_2_block_ram_r_5_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_6_0_inst : dff port map( d => n2493
                           , gclk => clk, rnot => n2365, q => 
                           load_n_store_RGB_Array_2_block_ram_r_6_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_6_1_inst : dff port map( d => n2494
                           , gclk => clk, rnot => n2366, q => 
                           load_n_store_RGB_Array_2_block_ram_r_6_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_6_2_inst : dff port map( d => n2495
                           , gclk => clk, rnot => n2367, q => 
                           load_n_store_RGB_Array_2_block_ram_r_6_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_6_3_inst : dff port map( d => n2496
                           , gclk => clk, rnot => n2368, q => 
                           load_n_store_RGB_Array_2_block_ram_r_6_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_6_4_inst : dff port map( d => n2497
                           , gclk => clk, rnot => n2369, q => 
                           load_n_store_RGB_Array_2_block_ram_r_6_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_6_5_inst : dff port map( d => n2498
                           , gclk => clk, rnot => n2370, q => 
                           load_n_store_RGB_Array_2_block_ram_r_6_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_6_6_inst : dff port map( d => n2499
                           , gclk => clk, rnot => n2371, q => 
                           load_n_store_RGB_Array_2_block_ram_r_6_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_6_7_inst : dff port map( d => n2500
                           , gclk => clk, rnot => n2372, q => 
                           load_n_store_RGB_Array_2_block_ram_r_6_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_7_0_inst : dff port map( d => n2501
                           , gclk => clk, rnot => n2373, q => 
                           load_n_store_RGB_Array_2_block_ram_r_7_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_7_1_inst : dff port map( d => n2502
                           , gclk => clk, rnot => n2374, q => 
                           load_n_store_RGB_Array_2_block_ram_r_7_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_7_2_inst : dff port map( d => n2503
                           , gclk => clk, rnot => n2375, q => 
                           load_n_store_RGB_Array_2_block_ram_r_7_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_7_3_inst : dff port map( d => n2504
                           , gclk => clk, rnot => n2376, q => 
                           load_n_store_RGB_Array_2_block_ram_r_7_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_7_4_inst : dff port map( d => n2505
                           , gclk => clk, rnot => n2377, q => 
                           load_n_store_RGB_Array_2_block_ram_r_7_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_7_5_inst : dff port map( d => n2506
                           , gclk => clk, rnot => n2378, q => 
                           load_n_store_RGB_Array_2_block_ram_r_7_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_7_6_inst : dff port map( d => n2507
                           , gclk => clk, rnot => n2379, q => 
                           load_n_store_RGB_Array_2_block_ram_r_7_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_7_7_inst : dff port map( d => n2508
                           , gclk => clk, rnot => n2380, q => 
                           load_n_store_RGB_Array_2_block_ram_r_7_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_8_0_inst : dff port map( d => n2509
                           , gclk => clk, rnot => n2381, q => 
                           load_n_store_RGB_Array_2_block_ram_r_8_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_8_1_inst : dff port map( d => n2510
                           , gclk => clk, rnot => n2382, q => 
                           load_n_store_RGB_Array_2_block_ram_r_8_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_8_2_inst : dff port map( d => n2511
                           , gclk => clk, rnot => n2383, q => 
                           load_n_store_RGB_Array_2_block_ram_r_8_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_8_3_inst : dff port map( d => n2512
                           , gclk => clk, rnot => n2384, q => 
                           load_n_store_RGB_Array_2_block_ram_r_8_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_8_4_inst : dff port map( d => n2513
                           , gclk => clk, rnot => n2385, q => 
                           load_n_store_RGB_Array_2_block_ram_r_8_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_8_5_inst : dff port map( d => n2514
                           , gclk => clk, rnot => n2386, q => 
                           load_n_store_RGB_Array_2_block_ram_r_8_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_8_6_inst : dff port map( d => n2515
                           , gclk => clk, rnot => n2387, q => 
                           load_n_store_RGB_Array_2_block_ram_r_8_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_8_7_inst : dff port map( d => n2516
                           , gclk => clk, rnot => n2388, q => 
                           load_n_store_RGB_Array_2_block_ram_r_8_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_9_0_inst : dff port map( d => n2517
                           , gclk => clk, rnot => n2389, q => 
                           load_n_store_RGB_Array_2_block_ram_r_9_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_9_1_inst : dff port map( d => n2518
                           , gclk => clk, rnot => n2390, q => 
                           load_n_store_RGB_Array_2_block_ram_r_9_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_9_2_inst : dff port map( d => n2519
                           , gclk => clk, rnot => n2391, q => 
                           load_n_store_RGB_Array_2_block_ram_r_9_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_9_3_inst : dff port map( d => n2520
                           , gclk => clk, rnot => n2392, q => 
                           load_n_store_RGB_Array_2_block_ram_r_9_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_9_4_inst : dff port map( d => n2521
                           , gclk => clk, rnot => n2393, q => 
                           load_n_store_RGB_Array_2_block_ram_r_9_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_9_5_inst : dff port map( d => n2522
                           , gclk => clk, rnot => n2394, q => 
                           load_n_store_RGB_Array_2_block_ram_r_9_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_9_6_inst : dff port map( d => n2523
                           , gclk => clk, rnot => n2395, q => 
                           load_n_store_RGB_Array_2_block_ram_r_9_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_9_7_inst : dff port map( d => n2524
                           , gclk => clk, rnot => n2396, q => 
                           load_n_store_RGB_Array_2_block_ram_r_9_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_10_0_inst : dff port map( d => 
                           n2525, gclk => clk, rnot => n2397, q => 
                           load_n_store_RGB_Array_2_block_ram_r_10_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_10_1_inst : dff port map( d => 
                           n2526, gclk => clk, rnot => n2398, q => 
                           load_n_store_RGB_Array_2_block_ram_r_10_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_10_2_inst : dff port map( d => 
                           n2527, gclk => clk, rnot => n2399, q => 
                           load_n_store_RGB_Array_2_block_ram_r_10_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_10_3_inst : dff port map( d => 
                           n2528, gclk => clk, rnot => n2400, q => 
                           load_n_store_RGB_Array_2_block_ram_r_10_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_10_4_inst : dff port map( d => 
                           n2529, gclk => clk, rnot => n2401, q => 
                           load_n_store_RGB_Array_2_block_ram_r_10_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_10_5_inst : dff port map( d => 
                           n2530, gclk => clk, rnot => n2402, q => 
                           load_n_store_RGB_Array_2_block_ram_r_10_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_10_6_inst : dff port map( d => 
                           n2531, gclk => clk, rnot => n2403, q => 
                           load_n_store_RGB_Array_2_block_ram_r_10_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_10_7_inst : dff port map( d => 
                           n2532, gclk => clk, rnot => n2404, q => 
                           load_n_store_RGB_Array_2_block_ram_r_10_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_11_0_inst : dff port map( d => 
                           n2533, gclk => clk, rnot => n2405, q => 
                           load_n_store_RGB_Array_2_block_ram_r_11_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_11_1_inst : dff port map( d => 
                           n2534, gclk => clk, rnot => n2406, q => 
                           load_n_store_RGB_Array_2_block_ram_r_11_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_11_2_inst : dff port map( d => 
                           n2535, gclk => clk, rnot => n2407, q => 
                           load_n_store_RGB_Array_2_block_ram_r_11_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_11_3_inst : dff port map( d => 
                           n2536, gclk => clk, rnot => n2408, q => 
                           load_n_store_RGB_Array_2_block_ram_r_11_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_11_4_inst : dff port map( d => 
                           n2537, gclk => clk, rnot => n2409, q => 
                           load_n_store_RGB_Array_2_block_ram_r_11_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_11_5_inst : dff port map( d => 
                           n2538, gclk => clk, rnot => n2410, q => 
                           load_n_store_RGB_Array_2_block_ram_r_11_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_11_6_inst : dff port map( d => 
                           n2539, gclk => clk, rnot => n2411, q => 
                           load_n_store_RGB_Array_2_block_ram_r_11_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_11_7_inst : dff port map( d => 
                           n2540, gclk => clk, rnot => n2412, q => 
                           load_n_store_RGB_Array_2_block_ram_r_11_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_12_0_inst : dff port map( d => 
                           n2541, gclk => clk, rnot => n2413, q => 
                           load_n_store_RGB_Array_2_block_ram_r_12_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_12_1_inst : dff port map( d => 
                           n2542, gclk => clk, rnot => n2414, q => 
                           load_n_store_RGB_Array_2_block_ram_r_12_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_12_2_inst : dff port map( d => 
                           n2543, gclk => clk, rnot => n2415, q => 
                           load_n_store_RGB_Array_2_block_ram_r_12_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_12_3_inst : dff port map( d => 
                           n2544, gclk => clk, rnot => n2416, q => 
                           load_n_store_RGB_Array_2_block_ram_r_12_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_12_4_inst : dff port map( d => 
                           n2545, gclk => clk, rnot => n2417, q => 
                           load_n_store_RGB_Array_2_block_ram_r_12_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_12_5_inst : dff port map( d => 
                           n2546, gclk => clk, rnot => n2418, q => 
                           load_n_store_RGB_Array_2_block_ram_r_12_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_12_6_inst : dff port map( d => 
                           n2547, gclk => clk, rnot => n2419, q => 
                           load_n_store_RGB_Array_2_block_ram_r_12_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_12_7_inst : dff port map( d => 
                           n2548, gclk => clk, rnot => n2420, q => 
                           load_n_store_RGB_Array_2_block_ram_r_12_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_13_0_inst : dff port map( d => 
                           n2549, gclk => clk, rnot => n2421, q => 
                           load_n_store_RGB_Array_2_block_ram_r_13_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_13_1_inst : dff port map( d => 
                           n2550, gclk => clk, rnot => n2422, q => 
                           load_n_store_RGB_Array_2_block_ram_r_13_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_13_2_inst : dff port map( d => 
                           n2551, gclk => clk, rnot => n2423, q => 
                           load_n_store_RGB_Array_2_block_ram_r_13_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_13_3_inst : dff port map( d => 
                           n2552, gclk => clk, rnot => n2424, q => 
                           load_n_store_RGB_Array_2_block_ram_r_13_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_13_4_inst : dff port map( d => 
                           n2553, gclk => clk, rnot => n2425, q => 
                           load_n_store_RGB_Array_2_block_ram_r_13_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_13_5_inst : dff port map( d => 
                           n2554, gclk => clk, rnot => n2426, q => 
                           load_n_store_RGB_Array_2_block_ram_r_13_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_13_6_inst : dff port map( d => 
                           n2555, gclk => clk, rnot => n2427, q => 
                           load_n_store_RGB_Array_2_block_ram_r_13_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_13_7_inst : dff port map( d => 
                           n2556, gclk => clk, rnot => n2428, q => 
                           load_n_store_RGB_Array_2_block_ram_r_13_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_14_0_inst : dff port map( d => 
                           n2557, gclk => clk, rnot => n2429, q => 
                           load_n_store_RGB_Array_2_block_ram_r_14_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_14_1_inst : dff port map( d => 
                           n2558, gclk => clk, rnot => n2430, q => 
                           load_n_store_RGB_Array_2_block_ram_r_14_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_14_2_inst : dff port map( d => 
                           n2559, gclk => clk, rnot => n2431, q => 
                           load_n_store_RGB_Array_2_block_ram_r_14_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_14_3_inst : dff port map( d => 
                           n2560, gclk => clk, rnot => n2432, q => 
                           load_n_store_RGB_Array_2_block_ram_r_14_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_14_4_inst : dff port map( d => 
                           n2561, gclk => clk, rnot => n2433, q => 
                           load_n_store_RGB_Array_2_block_ram_r_14_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_14_5_inst : dff port map( d => 
                           n2562, gclk => clk, rnot => n2434, q => 
                           load_n_store_RGB_Array_2_block_ram_r_14_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_14_6_inst : dff port map( d => 
                           n2563, gclk => clk, rnot => n2435, q => 
                           load_n_store_RGB_Array_2_block_ram_r_14_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_14_7_inst : dff port map( d => 
                           n2564, gclk => clk, rnot => n2436, q => 
                           load_n_store_RGB_Array_2_block_ram_r_14_7_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_15_0_inst : dff port map( d => 
                           n2565, gclk => clk, rnot => n2437, q => 
                           load_n_store_RGB_Array_2_block_ram_r_15_0_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_15_1_inst : dff port map( d => 
                           n2566, gclk => clk, rnot => n2438, q => 
                           load_n_store_RGB_Array_2_block_ram_r_15_1_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_15_2_inst : dff port map( d => 
                           n2567, gclk => clk, rnot => n2439, q => 
                           load_n_store_RGB_Array_2_block_ram_r_15_2_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_15_3_inst : dff port map( d => 
                           n2568, gclk => clk, rnot => n2440, q => 
                           load_n_store_RGB_Array_2_block_ram_r_15_3_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_15_4_inst : dff port map( d => 
                           n2569, gclk => clk, rnot => n2441, q => 
                           load_n_store_RGB_Array_2_block_ram_r_15_4_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_15_5_inst : dff port map( d => 
                           n2570, gclk => clk, rnot => n2442, q => 
                           load_n_store_RGB_Array_2_block_ram_r_15_5_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_15_6_inst : dff port map( d => 
                           n2571, gclk => clk, rnot => n2443, q => 
                           load_n_store_RGB_Array_2_block_ram_r_15_6_port);
   load_n_store_RGB_Array_2_block_ram_r_reg_15_7_inst : dff port map( d => 
                           n2572, gclk => clk, rnot => n2444, q => 
                           load_n_store_RGB_Array_2_block_ram_r_15_7_port);
   n2172 <= '1';
   n2171 <= '1';
   n2170 <= '1';
   n2169 <= '1';
   n2168 <= '1';
   n2167 <= '1';
   n2166 <= '1';
   n2165 <= '1';
   n2164 <= '1';
   n2163 <= '1';
   n2162 <= '1';
   n2161 <= '1';
   n2160 <= '1';
   n2159 <= '1';
   n2158 <= '1';
   n2157 <= '1';
   n2156 <= '1';
   n2155 <= '1';
   n2154 <= '1';
   n2153 <= '1';
   n2152 <= '1';
   n2151 <= '1';
   n2150 <= '1';
   n2149 <= '1';
   n2148 <= '1';
   n2147 <= '1';
   n2146 <= '1';
   n2145 <= '1';
   n2144 <= '1';
   n2143 <= '1';
   n2142 <= '1';
   n2141 <= '1';
   n2140 <= '1';
   n2139 <= '1';
   n2138 <= '1';
   n2137 <= '1';
   n2136 <= '1';
   n2135 <= '1';
   n2134 <= '1';
   n2133 <= '1';
   n2132 <= '1';
   n2131 <= '1';
   n2130 <= '1';
   n2129 <= '1';
   n2128 <= '1';
   n2127 <= '1';
   n2126 <= '1';
   n2125 <= '1';
   n2124 <= '1';
   n2123 <= '1';
   n2122 <= '1';
   n2121 <= '1';
   n2120 <= '1';
   n2119 <= '1';
   n2118 <= '1';
   n2117 <= '1';
   n2116 <= '1';
   n2115 <= '1';
   n2114 <= '1';
   n2113 <= '1';
   n2112 <= '1';
   n2111 <= '1';
   n2110 <= '1';
   n2109 <= '1';
   n2108 <= '1';
   n2107 <= '1';
   n2106 <= '1';
   n2105 <= '1';
   n2104 <= '1';
   n2103 <= '1';
   n2102 <= '1';
   n2101 <= '1';
   n2100 <= '1';
   n2099 <= '1';
   n2098 <= '1';
   n2097 <= '1';
   n2096 <= '1';
   n2095 <= '1';
   n2094 <= '1';
   n2093 <= '1';
   n2092 <= '1';
   n2091 <= '1';
   n2090 <= '1';
   n2089 <= '1';
   n2088 <= '1';
   n2087 <= '1';
   n2086 <= '1';
   n2085 <= '1';
   n2084 <= '1';
   n2083 <= '1';
   n2082 <= '1';
   n2081 <= '1';
   n2080 <= '1';
   n2079 <= '1';
   n2078 <= '1';
   n2077 <= '1';
   n2076 <= '1';
   n2075 <= '1';
   n2074 <= '1';
   n2073 <= '1';
   n2072 <= '1';
   n2071 <= '1';
   n2070 <= '1';
   n2069 <= '1';
   n2068 <= '1';
   n2067 <= '1';
   n2066 <= '1';
   n2065 <= '1';
   n2064 <= '1';
   n2063 <= '1';
   n2062 <= '1';
   n2061 <= '1';
   n2060 <= '1';
   n2059 <= '1';
   n2058 <= '1';
   n2057 <= '1';
   n2056 <= '1';
   n2055 <= '1';
   n2054 <= '1';
   n2053 <= '1';
   n2052 <= '1';
   n2051 <= '1';
   n2050 <= '1';
   n2049 <= '1';
   n2048 <= '1';
   n2047 <= '1';
   n2046 <= '1';
   n2045 <= '1';
   n2044 <= '1';
   n2043 <= '1';
   n2042 <= '1';
   n2041 <= '1';
   n2040 <= '1';
   n2039 <= '1';
   n2038 <= '1';
   n2037 <= '1';
   load_n_store_RGB_Array_1_data_out_o_reg_0_inst : dff port map( d => n2029, 
                           gclk => clk, rnot => n2037, q => 
                           load_n_store_lazy_out_1_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_0_0_inst : dff port map( d => n2173
                           , gclk => clk, rnot => n2038, q => 
                           load_n_store_RGB_Array_1_block_ram_r_0_0_port);
   load_n_store_RGB_Array_1_data_out_o_reg_1_inst : dff port map( d => n2030, 
                           gclk => clk, rnot => n2039, q => 
                           load_n_store_lazy_out_1_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_0_1_inst : dff port map( d => n2174
                           , gclk => clk, rnot => n2040, q => 
                           load_n_store_RGB_Array_1_block_ram_r_0_1_port);
   load_n_store_RGB_Array_1_data_out_o_reg_2_inst : dff port map( d => n2031, 
                           gclk => clk, rnot => n2041, q => 
                           load_n_store_lazy_out_1_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_0_2_inst : dff port map( d => n2175
                           , gclk => clk, rnot => n2042, q => 
                           load_n_store_RGB_Array_1_block_ram_r_0_2_port);
   load_n_store_RGB_Array_1_data_out_o_reg_3_inst : dff port map( d => n2032, 
                           gclk => clk, rnot => n2043, q => 
                           load_n_store_lazy_out_1_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_0_3_inst : dff port map( d => n2176
                           , gclk => clk, rnot => n2044, q => 
                           load_n_store_RGB_Array_1_block_ram_r_0_3_port);
   load_n_store_RGB_Array_1_data_out_o_reg_4_inst : dff port map( d => n2033, 
                           gclk => clk, rnot => n2045, q => 
                           load_n_store_lazy_out_1_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_0_4_inst : dff port map( d => n2177
                           , gclk => clk, rnot => n2046, q => 
                           load_n_store_RGB_Array_1_block_ram_r_0_4_port);
   load_n_store_RGB_Array_1_data_out_o_reg_5_inst : dff port map( d => n2034, 
                           gclk => clk, rnot => n2047, q => 
                           load_n_store_lazy_out_1_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_0_5_inst : dff port map( d => n2178
                           , gclk => clk, rnot => n2048, q => 
                           load_n_store_RGB_Array_1_block_ram_r_0_5_port);
   load_n_store_RGB_Array_1_data_out_o_reg_6_inst : dff port map( d => n2035, 
                           gclk => clk, rnot => n2049, q => 
                           load_n_store_lazy_out_1_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_0_6_inst : dff port map( d => n2179
                           , gclk => clk, rnot => n2050, q => 
                           load_n_store_RGB_Array_1_block_ram_r_0_6_port);
   load_n_store_RGB_Array_1_data_out_o_reg_7_inst : dff port map( d => n2036, 
                           gclk => clk, rnot => n2051, q => 
                           load_n_store_lazy_out_1_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_0_7_inst : dff port map( d => n2180
                           , gclk => clk, rnot => n2052, q => 
                           load_n_store_RGB_Array_1_block_ram_r_0_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_1_0_inst : dff port map( d => n2181
                           , gclk => clk, rnot => n2053, q => 
                           load_n_store_RGB_Array_1_block_ram_r_1_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_1_1_inst : dff port map( d => n2182
                           , gclk => clk, rnot => n2054, q => 
                           load_n_store_RGB_Array_1_block_ram_r_1_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_1_2_inst : dff port map( d => n2183
                           , gclk => clk, rnot => n2055, q => 
                           load_n_store_RGB_Array_1_block_ram_r_1_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_1_3_inst : dff port map( d => n2184
                           , gclk => clk, rnot => n2056, q => 
                           load_n_store_RGB_Array_1_block_ram_r_1_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_1_4_inst : dff port map( d => n2185
                           , gclk => clk, rnot => n2057, q => 
                           load_n_store_RGB_Array_1_block_ram_r_1_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_1_5_inst : dff port map( d => n2186
                           , gclk => clk, rnot => n2058, q => 
                           load_n_store_RGB_Array_1_block_ram_r_1_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_1_6_inst : dff port map( d => n2187
                           , gclk => clk, rnot => n2059, q => 
                           load_n_store_RGB_Array_1_block_ram_r_1_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_1_7_inst : dff port map( d => n2188
                           , gclk => clk, rnot => n2060, q => 
                           load_n_store_RGB_Array_1_block_ram_r_1_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_2_0_inst : dff port map( d => n2189
                           , gclk => clk, rnot => n2061, q => 
                           load_n_store_RGB_Array_1_block_ram_r_2_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_2_1_inst : dff port map( d => n2190
                           , gclk => clk, rnot => n2062, q => 
                           load_n_store_RGB_Array_1_block_ram_r_2_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_2_2_inst : dff port map( d => n2191
                           , gclk => clk, rnot => n2063, q => 
                           load_n_store_RGB_Array_1_block_ram_r_2_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_2_3_inst : dff port map( d => n2192
                           , gclk => clk, rnot => n2064, q => 
                           load_n_store_RGB_Array_1_block_ram_r_2_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_2_4_inst : dff port map( d => n2193
                           , gclk => clk, rnot => n2065, q => 
                           load_n_store_RGB_Array_1_block_ram_r_2_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_2_5_inst : dff port map( d => n2194
                           , gclk => clk, rnot => n2066, q => 
                           load_n_store_RGB_Array_1_block_ram_r_2_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_2_6_inst : dff port map( d => n2195
                           , gclk => clk, rnot => n2067, q => 
                           load_n_store_RGB_Array_1_block_ram_r_2_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_2_7_inst : dff port map( d => n2196
                           , gclk => clk, rnot => n2068, q => 
                           load_n_store_RGB_Array_1_block_ram_r_2_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_3_0_inst : dff port map( d => n2197
                           , gclk => clk, rnot => n2069, q => 
                           load_n_store_RGB_Array_1_block_ram_r_3_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_3_1_inst : dff port map( d => n2198
                           , gclk => clk, rnot => n2070, q => 
                           load_n_store_RGB_Array_1_block_ram_r_3_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_3_2_inst : dff port map( d => n2199
                           , gclk => clk, rnot => n2071, q => 
                           load_n_store_RGB_Array_1_block_ram_r_3_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_3_3_inst : dff port map( d => n2200
                           , gclk => clk, rnot => n2072, q => 
                           load_n_store_RGB_Array_1_block_ram_r_3_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_3_4_inst : dff port map( d => n2201
                           , gclk => clk, rnot => n2073, q => 
                           load_n_store_RGB_Array_1_block_ram_r_3_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_3_5_inst : dff port map( d => n2202
                           , gclk => clk, rnot => n2074, q => 
                           load_n_store_RGB_Array_1_block_ram_r_3_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_3_6_inst : dff port map( d => n2203
                           , gclk => clk, rnot => n2075, q => 
                           load_n_store_RGB_Array_1_block_ram_r_3_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_3_7_inst : dff port map( d => n2204
                           , gclk => clk, rnot => n2076, q => 
                           load_n_store_RGB_Array_1_block_ram_r_3_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_4_0_inst : dff port map( d => n2205
                           , gclk => clk, rnot => n2077, q => 
                           load_n_store_RGB_Array_1_block_ram_r_4_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_4_1_inst : dff port map( d => n2206
                           , gclk => clk, rnot => n2078, q => 
                           load_n_store_RGB_Array_1_block_ram_r_4_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_4_2_inst : dff port map( d => n2207
                           , gclk => clk, rnot => n2079, q => 
                           load_n_store_RGB_Array_1_block_ram_r_4_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_4_3_inst : dff port map( d => n2208
                           , gclk => clk, rnot => n2080, q => 
                           load_n_store_RGB_Array_1_block_ram_r_4_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_4_4_inst : dff port map( d => n2209
                           , gclk => clk, rnot => n2081, q => 
                           load_n_store_RGB_Array_1_block_ram_r_4_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_4_5_inst : dff port map( d => n2210
                           , gclk => clk, rnot => n2082, q => 
                           load_n_store_RGB_Array_1_block_ram_r_4_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_4_6_inst : dff port map( d => n2211
                           , gclk => clk, rnot => n2083, q => 
                           load_n_store_RGB_Array_1_block_ram_r_4_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_4_7_inst : dff port map( d => n2212
                           , gclk => clk, rnot => n2084, q => 
                           load_n_store_RGB_Array_1_block_ram_r_4_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_5_0_inst : dff port map( d => n2213
                           , gclk => clk, rnot => n2085, q => 
                           load_n_store_RGB_Array_1_block_ram_r_5_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_5_1_inst : dff port map( d => n2214
                           , gclk => clk, rnot => n2086, q => 
                           load_n_store_RGB_Array_1_block_ram_r_5_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_5_2_inst : dff port map( d => n2215
                           , gclk => clk, rnot => n2087, q => 
                           load_n_store_RGB_Array_1_block_ram_r_5_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_5_3_inst : dff port map( d => n2216
                           , gclk => clk, rnot => n2088, q => 
                           load_n_store_RGB_Array_1_block_ram_r_5_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_5_4_inst : dff port map( d => n2217
                           , gclk => clk, rnot => n2089, q => 
                           load_n_store_RGB_Array_1_block_ram_r_5_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_5_5_inst : dff port map( d => n2218
                           , gclk => clk, rnot => n2090, q => 
                           load_n_store_RGB_Array_1_block_ram_r_5_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_5_6_inst : dff port map( d => n2219
                           , gclk => clk, rnot => n2091, q => 
                           load_n_store_RGB_Array_1_block_ram_r_5_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_5_7_inst : dff port map( d => n2220
                           , gclk => clk, rnot => n2092, q => 
                           load_n_store_RGB_Array_1_block_ram_r_5_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_6_0_inst : dff port map( d => n2221
                           , gclk => clk, rnot => n2093, q => 
                           load_n_store_RGB_Array_1_block_ram_r_6_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_6_1_inst : dff port map( d => n2222
                           , gclk => clk, rnot => n2094, q => 
                           load_n_store_RGB_Array_1_block_ram_r_6_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_6_2_inst : dff port map( d => n2223
                           , gclk => clk, rnot => n2095, q => 
                           load_n_store_RGB_Array_1_block_ram_r_6_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_6_3_inst : dff port map( d => n2224
                           , gclk => clk, rnot => n2096, q => 
                           load_n_store_RGB_Array_1_block_ram_r_6_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_6_4_inst : dff port map( d => n2225
                           , gclk => clk, rnot => n2097, q => 
                           load_n_store_RGB_Array_1_block_ram_r_6_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_6_5_inst : dff port map( d => n2226
                           , gclk => clk, rnot => n2098, q => 
                           load_n_store_RGB_Array_1_block_ram_r_6_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_6_6_inst : dff port map( d => n2227
                           , gclk => clk, rnot => n2099, q => 
                           load_n_store_RGB_Array_1_block_ram_r_6_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_6_7_inst : dff port map( d => n2228
                           , gclk => clk, rnot => n2100, q => 
                           load_n_store_RGB_Array_1_block_ram_r_6_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_7_0_inst : dff port map( d => n2229
                           , gclk => clk, rnot => n2101, q => 
                           load_n_store_RGB_Array_1_block_ram_r_7_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_7_1_inst : dff port map( d => n2230
                           , gclk => clk, rnot => n2102, q => 
                           load_n_store_RGB_Array_1_block_ram_r_7_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_7_2_inst : dff port map( d => n2231
                           , gclk => clk, rnot => n2103, q => 
                           load_n_store_RGB_Array_1_block_ram_r_7_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_7_3_inst : dff port map( d => n2232
                           , gclk => clk, rnot => n2104, q => 
                           load_n_store_RGB_Array_1_block_ram_r_7_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_7_4_inst : dff port map( d => n2233
                           , gclk => clk, rnot => n2105, q => 
                           load_n_store_RGB_Array_1_block_ram_r_7_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_7_5_inst : dff port map( d => n2234
                           , gclk => clk, rnot => n2106, q => 
                           load_n_store_RGB_Array_1_block_ram_r_7_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_7_6_inst : dff port map( d => n2235
                           , gclk => clk, rnot => n2107, q => 
                           load_n_store_RGB_Array_1_block_ram_r_7_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_7_7_inst : dff port map( d => n2236
                           , gclk => clk, rnot => n2108, q => 
                           load_n_store_RGB_Array_1_block_ram_r_7_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_8_0_inst : dff port map( d => n2237
                           , gclk => clk, rnot => n2109, q => 
                           load_n_store_RGB_Array_1_block_ram_r_8_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_8_1_inst : dff port map( d => n2238
                           , gclk => clk, rnot => n2110, q => 
                           load_n_store_RGB_Array_1_block_ram_r_8_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_8_2_inst : dff port map( d => n2239
                           , gclk => clk, rnot => n2111, q => 
                           load_n_store_RGB_Array_1_block_ram_r_8_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_8_3_inst : dff port map( d => n2240
                           , gclk => clk, rnot => n2112, q => 
                           load_n_store_RGB_Array_1_block_ram_r_8_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_8_4_inst : dff port map( d => n2241
                           , gclk => clk, rnot => n2113, q => 
                           load_n_store_RGB_Array_1_block_ram_r_8_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_8_5_inst : dff port map( d => n2242
                           , gclk => clk, rnot => n2114, q => 
                           load_n_store_RGB_Array_1_block_ram_r_8_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_8_6_inst : dff port map( d => n2243
                           , gclk => clk, rnot => n2115, q => 
                           load_n_store_RGB_Array_1_block_ram_r_8_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_8_7_inst : dff port map( d => n2244
                           , gclk => clk, rnot => n2116, q => 
                           load_n_store_RGB_Array_1_block_ram_r_8_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_9_0_inst : dff port map( d => n2245
                           , gclk => clk, rnot => n2117, q => 
                           load_n_store_RGB_Array_1_block_ram_r_9_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_9_1_inst : dff port map( d => n2246
                           , gclk => clk, rnot => n2118, q => 
                           load_n_store_RGB_Array_1_block_ram_r_9_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_9_2_inst : dff port map( d => n2247
                           , gclk => clk, rnot => n2119, q => 
                           load_n_store_RGB_Array_1_block_ram_r_9_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_9_3_inst : dff port map( d => n2248
                           , gclk => clk, rnot => n2120, q => 
                           load_n_store_RGB_Array_1_block_ram_r_9_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_9_4_inst : dff port map( d => n2249
                           , gclk => clk, rnot => n2121, q => 
                           load_n_store_RGB_Array_1_block_ram_r_9_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_9_5_inst : dff port map( d => n2250
                           , gclk => clk, rnot => n2122, q => 
                           load_n_store_RGB_Array_1_block_ram_r_9_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_9_6_inst : dff port map( d => n2251
                           , gclk => clk, rnot => n2123, q => 
                           load_n_store_RGB_Array_1_block_ram_r_9_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_9_7_inst : dff port map( d => n2252
                           , gclk => clk, rnot => n2124, q => 
                           load_n_store_RGB_Array_1_block_ram_r_9_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_10_0_inst : dff port map( d => 
                           n2253, gclk => clk, rnot => n2125, q => 
                           load_n_store_RGB_Array_1_block_ram_r_10_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_10_1_inst : dff port map( d => 
                           n2254, gclk => clk, rnot => n2126, q => 
                           load_n_store_RGB_Array_1_block_ram_r_10_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_10_2_inst : dff port map( d => 
                           n2255, gclk => clk, rnot => n2127, q => 
                           load_n_store_RGB_Array_1_block_ram_r_10_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_10_3_inst : dff port map( d => 
                           n2256, gclk => clk, rnot => n2128, q => 
                           load_n_store_RGB_Array_1_block_ram_r_10_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_10_4_inst : dff port map( d => 
                           n2257, gclk => clk, rnot => n2129, q => 
                           load_n_store_RGB_Array_1_block_ram_r_10_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_10_5_inst : dff port map( d => 
                           n2258, gclk => clk, rnot => n2130, q => 
                           load_n_store_RGB_Array_1_block_ram_r_10_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_10_6_inst : dff port map( d => 
                           n2259, gclk => clk, rnot => n2131, q => 
                           load_n_store_RGB_Array_1_block_ram_r_10_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_10_7_inst : dff port map( d => 
                           n2260, gclk => clk, rnot => n2132, q => 
                           load_n_store_RGB_Array_1_block_ram_r_10_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_11_0_inst : dff port map( d => 
                           n2261, gclk => clk, rnot => n2133, q => 
                           load_n_store_RGB_Array_1_block_ram_r_11_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_11_1_inst : dff port map( d => 
                           n2262, gclk => clk, rnot => n2134, q => 
                           load_n_store_RGB_Array_1_block_ram_r_11_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_11_2_inst : dff port map( d => 
                           n2263, gclk => clk, rnot => n2135, q => 
                           load_n_store_RGB_Array_1_block_ram_r_11_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_11_3_inst : dff port map( d => 
                           n2264, gclk => clk, rnot => n2136, q => 
                           load_n_store_RGB_Array_1_block_ram_r_11_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_11_4_inst : dff port map( d => 
                           n2265, gclk => clk, rnot => n2137, q => 
                           load_n_store_RGB_Array_1_block_ram_r_11_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_11_5_inst : dff port map( d => 
                           n2266, gclk => clk, rnot => n2138, q => 
                           load_n_store_RGB_Array_1_block_ram_r_11_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_11_6_inst : dff port map( d => 
                           n2267, gclk => clk, rnot => n2139, q => 
                           load_n_store_RGB_Array_1_block_ram_r_11_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_11_7_inst : dff port map( d => 
                           n2268, gclk => clk, rnot => n2140, q => 
                           load_n_store_RGB_Array_1_block_ram_r_11_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_12_0_inst : dff port map( d => 
                           n2269, gclk => clk, rnot => n2141, q => 
                           load_n_store_RGB_Array_1_block_ram_r_12_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_12_1_inst : dff port map( d => 
                           n2270, gclk => clk, rnot => n2142, q => 
                           load_n_store_RGB_Array_1_block_ram_r_12_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_12_2_inst : dff port map( d => 
                           n2271, gclk => clk, rnot => n2143, q => 
                           load_n_store_RGB_Array_1_block_ram_r_12_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_12_3_inst : dff port map( d => 
                           n2272, gclk => clk, rnot => n2144, q => 
                           load_n_store_RGB_Array_1_block_ram_r_12_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_12_4_inst : dff port map( d => 
                           n2273, gclk => clk, rnot => n2145, q => 
                           load_n_store_RGB_Array_1_block_ram_r_12_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_12_5_inst : dff port map( d => 
                           n2274, gclk => clk, rnot => n2146, q => 
                           load_n_store_RGB_Array_1_block_ram_r_12_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_12_6_inst : dff port map( d => 
                           n2275, gclk => clk, rnot => n2147, q => 
                           load_n_store_RGB_Array_1_block_ram_r_12_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_12_7_inst : dff port map( d => 
                           n2276, gclk => clk, rnot => n2148, q => 
                           load_n_store_RGB_Array_1_block_ram_r_12_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_13_0_inst : dff port map( d => 
                           n2277, gclk => clk, rnot => n2149, q => 
                           load_n_store_RGB_Array_1_block_ram_r_13_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_13_1_inst : dff port map( d => 
                           n2278, gclk => clk, rnot => n2150, q => 
                           load_n_store_RGB_Array_1_block_ram_r_13_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_13_2_inst : dff port map( d => 
                           n2279, gclk => clk, rnot => n2151, q => 
                           load_n_store_RGB_Array_1_block_ram_r_13_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_13_3_inst : dff port map( d => 
                           n2280, gclk => clk, rnot => n2152, q => 
                           load_n_store_RGB_Array_1_block_ram_r_13_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_13_4_inst : dff port map( d => 
                           n2281, gclk => clk, rnot => n2153, q => 
                           load_n_store_RGB_Array_1_block_ram_r_13_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_13_5_inst : dff port map( d => 
                           n2282, gclk => clk, rnot => n2154, q => 
                           load_n_store_RGB_Array_1_block_ram_r_13_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_13_6_inst : dff port map( d => 
                           n2283, gclk => clk, rnot => n2155, q => 
                           load_n_store_RGB_Array_1_block_ram_r_13_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_13_7_inst : dff port map( d => 
                           n2284, gclk => clk, rnot => n2156, q => 
                           load_n_store_RGB_Array_1_block_ram_r_13_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_14_0_inst : dff port map( d => 
                           n2285, gclk => clk, rnot => n2157, q => 
                           load_n_store_RGB_Array_1_block_ram_r_14_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_14_1_inst : dff port map( d => 
                           n2286, gclk => clk, rnot => n2158, q => 
                           load_n_store_RGB_Array_1_block_ram_r_14_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_14_2_inst : dff port map( d => 
                           n2287, gclk => clk, rnot => n2159, q => 
                           load_n_store_RGB_Array_1_block_ram_r_14_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_14_3_inst : dff port map( d => 
                           n2288, gclk => clk, rnot => n2160, q => 
                           load_n_store_RGB_Array_1_block_ram_r_14_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_14_4_inst : dff port map( d => 
                           n2289, gclk => clk, rnot => n2161, q => 
                           load_n_store_RGB_Array_1_block_ram_r_14_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_14_5_inst : dff port map( d => 
                           n2290, gclk => clk, rnot => n2162, q => 
                           load_n_store_RGB_Array_1_block_ram_r_14_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_14_6_inst : dff port map( d => 
                           n2291, gclk => clk, rnot => n2163, q => 
                           load_n_store_RGB_Array_1_block_ram_r_14_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_14_7_inst : dff port map( d => 
                           n2292, gclk => clk, rnot => n2164, q => 
                           load_n_store_RGB_Array_1_block_ram_r_14_7_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_15_0_inst : dff port map( d => 
                           n2293, gclk => clk, rnot => n2165, q => 
                           load_n_store_RGB_Array_1_block_ram_r_15_0_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_15_1_inst : dff port map( d => 
                           n2294, gclk => clk, rnot => n2166, q => 
                           load_n_store_RGB_Array_1_block_ram_r_15_1_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_15_2_inst : dff port map( d => 
                           n2295, gclk => clk, rnot => n2167, q => 
                           load_n_store_RGB_Array_1_block_ram_r_15_2_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_15_3_inst : dff port map( d => 
                           n2296, gclk => clk, rnot => n2168, q => 
                           load_n_store_RGB_Array_1_block_ram_r_15_3_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_15_4_inst : dff port map( d => 
                           n2297, gclk => clk, rnot => n2169, q => 
                           load_n_store_RGB_Array_1_block_ram_r_15_4_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_15_5_inst : dff port map( d => 
                           n2298, gclk => clk, rnot => n2170, q => 
                           load_n_store_RGB_Array_1_block_ram_r_15_5_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_15_6_inst : dff port map( d => 
                           n2299, gclk => clk, rnot => n2171, q => 
                           load_n_store_RGB_Array_1_block_ram_r_15_6_port);
   load_n_store_RGB_Array_1_block_ram_r_reg_15_7_inst : dff port map( d => 
                           n2300, gclk => clk, rnot => n2172, q => 
                           load_n_store_RGB_Array_1_block_ram_r_15_7_port);
   U1 : oai22 port map( a => n1, b => n2, c => n3, d => n4, outb => 
                           registers_n286);
   U2 : nor2 port map( a => n5, b => n3, outb => n2);
   U3 : oai22 port map( a => n1, b => n6, c => n7, d => n8, outb => 
                           registers_n285);
   U4 : nor2 port map( a => n1, b => registers_s_delay_0_port, outb => n7);
   U5 : inv port map( inb => n4, outb => n1);
   U6 : oai12 port map( b => n9, c => n10, a => n11, outb => n4);
   U7 : nand3 port map( a => n11, b => n12, c => n13, outb => registers_n284);
   U8 : oai22 port map( a => n14, b => n15, c => n16, d => n17, outb => 
                           registers_n283);
   U9 : aoi12 port map( b => n18, c => n6, a => n19, outb => n16);
   U10 : oai22 port map( a => n20, b => n21, c => n22, d => n17, outb => 
                           registers_n282);
   U11 : oai12 port map( b => registers_reg_col_inc_0_port, c => n15, a => n23,
                           outb => registers_n281);
   U12 : nand3 port map( a => n18, b => n6, c => registers_reg_col_inc_0_port, 
                           outb => n23);
   U13 : inv port map( inb => n19, outb => n15);
   U14 : oai22 port map( a => n24, b => n21, c => n22, d => n14, outb => 
                           registers_n280);
   U15 : oai22 port map( a => n25, b => n26, c => n27, d => n28, outb => 
                           registers_n279);
   U16 : inv port map( inb => n29, outb => n27);
   U17 : nand2 port map( a => n30, b => n31, outb => n29);
   U18 : oai22 port map( a => n32, b => n30, c => registers_reg_cd_0_port, d =>
                           n26, outb => registers_n278);
   U19 : oai12 port map( b => n31, c => n33, a => n34, outb => registers_n277);
   U20 : inv port map( inb => n35, outb => n34);
   U21 : oai22 port map( a => n36, b => n26, c => n30, d => n37, outb => n35);
   U22 : nand2 port map( a => n38, b => n30, outb => n26);
   U23 : nand2 port map( a => n39, b => n11, outb => n30);
   U24 : inv port map( inb => n38, outb => n31);
   U25 : nor2 port map( a => n6, b => n40, outb => n38);
   U26 : oai12 port map( b => n41, c => n42, a => n43, outb => registers_n276);
   U27 : nand4 port map( a => n5, b => n44, c => registers_reg_row_0_port, d =>
                           n42, outb => n43);
   U28 : aoi12 port map( b => n5, c => n45, a => n39, outb => n41);
   U29 : inv port map( inb => n44, outb => n39);
   U30 : oai22 port map( a => n46, b => n21, c => n22, d => n42, outb => 
                           registers_n275);
   U31 : inv port map( inb => registers_reg_row_1_port, outb => n42);
   U32 : oai12 port map( b => n44, c => n45, a => n47, outb => registers_n274);
   U33 : nand3 port map( a => n5, b => n44, c => n45, outb => n47);
   U34 : oai12 port map( b => n48, c => n11, a => n18, outb => n44);
   U35 : inv port map( inb => n49, outb => n18);
   U36 : nand2 port map( a => n50, b => n51, outb => n11);
   U37 : oai22 port map( a => n52, b => n21, c => n22, d => n45, outb => 
                           registers_n273);
   U38 : inv port map( inb => registers_reg_row_0_port, outb => n45);
   U39 : inv port map( inb => n22, outb => n21);
   U40 : nor2 port map( a => n49, b => n50, outb => n22);
   U41 : nand3 port map( a => n53, b => n54, c => n12, outb => registers_n272);
   U42 : nand3 port map( a => n55, b => n56, c => mem_reg_f, outb => n12);
   U43 : nand2 port map( a => n55, b => n57, outb => n54);
   U44 : nand4 port map( a => n58, b => n6, c => reg_hub_f, d => n10, outb => 
                           n53);
   U45 : oai22 port map( a => n59, b => n60, c => n50, d => n61, outb => 
                           registers_n271);
   U46 : oai12 port map( b => mem_out_b0_7_port, c => n48, a => n62, outb => 
                           n60);
   U47 : aoi22 port map( a => registers_reg_cd_2_port, b => n63, c => n64, d =>
                           n28, outb => n62);
   U48 : inv port map( inb => n65, outb => n64);
   U49 : nor2 port map( a => n66, b => n67, outb => n65);
   U50 : oai22 port map( a => n25, b => mem_out_b0_3_port, c => n68, d => 
                           mem_out_b0_0_port, outb => n67);
   U51 : oai22 port map( a => n33, b => mem_out_b0_2_port, c => n36, d => 
                           mem_out_b0_1_port, outb => n66);
   U52 : oai12 port map( b => mem_out_b0_5_port, c => n36, a => n69, outb => 
                           n63);
   U53 : inv port map( inb => n70, outb => n69);
   U54 : oai22 port map( a => n33, b => mem_out_b0_6_port, c => n68, d => 
                           mem_out_b0_4_port, outb => n70);
   U55 : oai22 port map( a => n10, b => n61, c => n55, d => n71, outb => 
                           registers_n270);
   U56 : oai22 port map( a => n59, b => n61, c => n50, d => n72, outb => 
                           registers_n269);
   U57 : inv port map( inb => registers_s_mem_sipo_b0_7_port, outb => n61);
   U58 : inv port map( inb => n73, outb => registers_n268);
   U59 : aoi22 port map( a => n55, b => registers_s_mem_sipo_b0_6_port, c => 
                           n10, d => mem_sipo_b0_6_port, outb => n73);
   U60 : oai22 port map( a => n59, b => n72, c => n50, d => n74, outb => 
                           registers_n267);
   U61 : inv port map( inb => registers_s_mem_sipo_b0_6_port, outb => n72);
   U62 : inv port map( inb => n75, outb => registers_n266);
   U63 : aoi22 port map( a => n55, b => registers_s_mem_sipo_b0_5_port, c => 
                           n10, d => mem_sipo_b0_5_port, outb => n75);
   U64 : oai22 port map( a => n59, b => n74, c => n50, d => n76, outb => 
                           registers_n265);
   U65 : inv port map( inb => registers_s_mem_sipo_b0_5_port, outb => n74);
   U66 : inv port map( inb => n77, outb => registers_n264);
   U67 : aoi22 port map( a => n55, b => registers_s_mem_sipo_b0_4_port, c => 
                           n10, d => mem_sipo_b0_4_port, outb => n77);
   U68 : oai22 port map( a => n59, b => n76, c => n50, d => n78, outb => 
                           registers_n263);
   U69 : inv port map( inb => registers_s_mem_sipo_b0_4_port, outb => n76);
   U70 : inv port map( inb => n79, outb => registers_n262);
   U71 : aoi22 port map( a => n55, b => registers_s_mem_sipo_b0_3_port, c => 
                           n10, d => mem_sipo_b0_3_port, outb => n79);
   U72 : oai22 port map( a => n59, b => n78, c => n50, d => n80, outb => 
                           registers_n261);
   U73 : inv port map( inb => registers_s_mem_sipo_b0_3_port, outb => n78);
   U74 : inv port map( inb => n81, outb => registers_n260);
   U75 : aoi22 port map( a => n55, b => registers_s_mem_sipo_b0_2_port, c => 
                           n10, d => mem_sipo_b0_2_port, outb => n81);
   U76 : oai22 port map( a => n59, b => n80, c => n50, d => n82, outb => 
                           registers_n259);
   U77 : inv port map( inb => registers_s_mem_sipo_b0_2_port, outb => n80);
   U78 : oai22 port map( a => n10, b => n82, c => n55, d => n83, outb => 
                           registers_n258);
   U79 : inv port map( inb => mem_sipo_b0_1_port, outb => n83);
   U80 : inv port map( inb => registers_s_mem_sipo_b0_1_port, outb => n82);
   U81 : inv port map( inb => n84, outb => registers_n257);
   U82 : aoi22 port map( a => n50, b => registers_s_mem_sipo_b0_1_port, c => 
                           n59, d => registers_s_mem_sipo_b0_0_port, outb => 
                           n84);
   U83 : inv port map( inb => n85, outb => registers_n256);
   U84 : aoi22 port map( a => n55, b => registers_s_mem_sipo_b0_0_port, c => 
                           n10, d => mem_sipo_b0_0_port, outb => n85);
   U85 : oai22 port map( a => n59, b => n86, c => n50, d => n87, outb => 
                           registers_n255);
   U86 : oai12 port map( b => mem_out_r0_7_port, c => n48, a => n88, outb => 
                           n86);
   U87 : aoi22 port map( a => registers_reg_cd_2_port, b => n89, c => n90, d =>
                           n28, outb => n88);
   U88 : inv port map( inb => n91, outb => n90);
   U89 : nor2 port map( a => n92, b => n93, outb => n91);
   U90 : oai22 port map( a => n25, b => mem_out_r0_3_port, c => n68, d => 
                           mem_out_r0_0_port, outb => n93);
   U91 : oai22 port map( a => n33, b => mem_out_r0_2_port, c => n36, d => 
                           mem_out_r0_1_port, outb => n92);
   U92 : oai12 port map( b => mem_out_r0_5_port, c => n36, a => n94, outb => 
                           n89);
   U93 : inv port map( inb => n95, outb => n94);
   U94 : oai22 port map( a => n33, b => mem_out_r0_6_port, c => n68, d => 
                           mem_out_r0_4_port, outb => n95);
   U95 : oai22 port map( a => n59, b => n87, c => n50, d => n96, outb => 
                           registers_n254);
   U96 : oai22 port map( a => n59, b => n96, c => n50, d => n97, outb => 
                           registers_n253);
   U97 : inv port map( inb => registers_s_mem_sipo_r0_6_port, outb => n96);
   U98 : oai22 port map( a => n59, b => n97, c => n50, d => n98, outb => 
                           registers_n252);
   U99 : inv port map( inb => registers_s_mem_sipo_r0_5_port, outb => n97);
   U100 : oai22 port map( a => n59, b => n98, c => n50, d => n99, outb => 
                           registers_n251);
   U101 : inv port map( inb => registers_s_mem_sipo_r0_4_port, outb => n98);
   U102 : oai22 port map( a => n59, b => n99, c => n50, d => n100, outb => 
                           registers_n250);
   U103 : inv port map( inb => registers_s_mem_sipo_r0_3_port, outb => n99);
   U104 : oai22 port map( a => n59, b => n100, c => n50, d => n101, outb => 
                           registers_n249);
   U105 : inv port map( inb => registers_s_mem_sipo_r0_2_port, outb => n100);
   U106 : inv port map( inb => n102, outb => registers_n248);
   U107 : aoi22 port map( a => n50, b => registers_s_mem_sipo_r0_1_port, c => 
                           n59, d => registers_s_mem_sipo_r0_0_port, outb => 
                           n102);
   U108 : oai22 port map( a => n59, b => n103, c => n50, d => n104, outb => 
                           registers_n247);
   U109 : oai12 port map( b => mem_out_g0_7_port, c => n48, a => n105, outb => 
                           n103);
   U110 : aoi22 port map( a => registers_reg_cd_2_port, b => n106, c => n107, d
                           => n28, outb => n105);
   U111 : inv port map( inb => n108, outb => n107);
   U112 : nor2 port map( a => n109, b => n110, outb => n108);
   U113 : oai22 port map( a => n25, b => mem_out_g0_3_port, c => n68, d => 
                           mem_out_g0_0_port, outb => n110);
   U114 : oai22 port map( a => n33, b => mem_out_g0_2_port, c => n36, d => 
                           mem_out_g0_1_port, outb => n109);
   U115 : oai12 port map( b => mem_out_g0_5_port, c => n36, a => n111, outb => 
                           n106);
   U116 : inv port map( inb => n112, outb => n111);
   U117 : oai22 port map( a => n33, b => mem_out_g0_6_port, c => n68, d => 
                           mem_out_g0_4_port, outb => n112);
   U118 : nand2 port map( a => n37, b => n32, outb => n68);
   U119 : nand2 port map( a => registers_reg_cd_1_port, b => n32, outb => n33);
   U120 : inv port map( inb => registers_reg_cd_0_port, outb => n32);
   U121 : nand2 port map( a => registers_reg_cd_0_port, b => n37, outb => n36);
   U122 : inv port map( inb => registers_reg_cd_1_port, outb => n37);
   U123 : inv port map( inb => n40, outb => n48);
   U124 : nor2 port map( a => n28, b => n25, outb => n40);
   U125 : nand2 port map( a => registers_reg_cd_1_port, b => 
                           registers_reg_cd_0_port, outb => n25);
   U126 : inv port map( inb => registers_reg_cd_2_port, outb => n28);
   U127 : oai22 port map( a => n59, b => n104, c => n50, d => n113, outb => 
                           registers_n246);
   U128 : oai22 port map( a => n59, b => n113, c => n50, d => n114, outb => 
                           registers_n245);
   U129 : inv port map( inb => registers_s_mem_sipo_g0_6_port, outb => n113);
   U130 : oai22 port map( a => n59, b => n114, c => n50, d => n115, outb => 
                           registers_n244);
   U131 : inv port map( inb => registers_s_mem_sipo_g0_5_port, outb => n114);
   U132 : oai22 port map( a => n59, b => n115, c => n50, d => n116, outb => 
                           registers_n243);
   U133 : inv port map( inb => registers_s_mem_sipo_g0_4_port, outb => n115);
   U134 : oai22 port map( a => n59, b => n116, c => n50, d => n117, outb => 
                           registers_n242);
   U135 : inv port map( inb => registers_s_mem_sipo_g0_3_port, outb => n116);
   U136 : oai22 port map( a => n59, b => n117, c => n50, d => n118, outb => 
                           registers_n241);
   U137 : inv port map( inb => registers_s_mem_sipo_g0_2_port, outb => n117);
   U138 : inv port map( inb => n119, outb => registers_n240);
   U139 : aoi22 port map( a => n50, b => registers_s_mem_sipo_g0_1_port, c => 
                           n59, d => registers_s_mem_sipo_g0_0_port, outb => 
                           n119);
   U140 : oai22 port map( a => n10, b => n87, c => n55, d => n120, outb => 
                           registers_n239);
   U141 : inv port map( inb => registers_s_mem_sipo_r0_7_port, outb => n87);
   U142 : inv port map( inb => n121, outb => registers_n238);
   U143 : aoi22 port map( a => n55, b => registers_s_mem_sipo_r0_6_port, c => 
                           n10, d => mem_sipo_r0_6_port, outb => n121);
   U144 : inv port map( inb => n122, outb => registers_n237);
   U145 : aoi22 port map( a => n55, b => registers_s_mem_sipo_r0_5_port, c => 
                           n10, d => mem_sipo_r0_5_port, outb => n122);
   U146 : inv port map( inb => n123, outb => registers_n236);
   U147 : aoi22 port map( a => n55, b => registers_s_mem_sipo_r0_4_port, c => 
                           n10, d => mem_sipo_r0_4_port, outb => n123);
   U148 : inv port map( inb => n124, outb => registers_n235);
   U149 : aoi22 port map( a => n55, b => registers_s_mem_sipo_r0_3_port, c => 
                           n10, d => mem_sipo_r0_3_port, outb => n124);
   U150 : inv port map( inb => n125, outb => registers_n234);
   U151 : aoi22 port map( a => n55, b => registers_s_mem_sipo_r0_2_port, c => 
                           n10, d => mem_sipo_r0_2_port, outb => n125);
   U152 : oai22 port map( a => n10, b => n101, c => n55, d => n126, outb => 
                           registers_n233);
   U153 : inv port map( inb => mem_sipo_r0_1_port, outb => n126);
   U154 : inv port map( inb => registers_s_mem_sipo_r0_1_port, outb => n101);
   U155 : inv port map( inb => n127, outb => registers_n232);
   U156 : aoi22 port map( a => n55, b => registers_s_mem_sipo_r0_0_port, c => 
                           n10, d => mem_sipo_r0_0_port, outb => n127);
   U157 : oai22 port map( a => n10, b => n104, c => n55, d => n128, outb => 
                           registers_n231);
   U158 : inv port map( inb => registers_s_mem_sipo_g0_7_port, outb => n104);
   U159 : inv port map( inb => n129, outb => registers_n230);
   U160 : aoi22 port map( a => n55, b => registers_s_mem_sipo_g0_6_port, c => 
                           n10, d => mem_sipo_g0_6_port, outb => n129);
   U161 : inv port map( inb => n130, outb => registers_n229);
   U162 : aoi22 port map( a => n55, b => registers_s_mem_sipo_g0_5_port, c => 
                           n10, d => mem_sipo_g0_5_port, outb => n130);
   U163 : inv port map( inb => n131, outb => registers_n228);
   U164 : aoi22 port map( a => n55, b => registers_s_mem_sipo_g0_4_port, c => 
                           n10, d => mem_sipo_g0_4_port, outb => n131);
   U165 : inv port map( inb => n132, outb => registers_n227);
   U166 : aoi22 port map( a => n55, b => registers_s_mem_sipo_g0_3_port, c => 
                           n10, d => mem_sipo_g0_3_port, outb => n132);
   U167 : inv port map( inb => n133, outb => registers_n226);
   U168 : aoi22 port map( a => n55, b => registers_s_mem_sipo_g0_2_port, c => 
                           n10, d => mem_sipo_g0_2_port, outb => n133);
   U169 : oai22 port map( a => n10, b => n118, c => n55, d => n134, outb => 
                           registers_n225);
   U170 : inv port map( inb => mem_sipo_g0_1_port, outb => n134);
   U171 : inv port map( inb => registers_s_mem_sipo_g0_1_port, outb => n118);
   U172 : inv port map( inb => n135, outb => registers_n224);
   U173 : aoi22 port map( a => n55, b => registers_s_mem_sipo_g0_0_port, c => 
                           n10, d => mem_sipo_g0_0_port, outb => n135);
   U174 : oai22 port map( a => n136, b => n137, c => n138, d => n139, outb => 
                           n1894);
   U175 : inv port map( inb => n137, outb => n138);
   U176 : nand2 port map( a => n140, b => n141, outb => n137);
   U177 : inv port map( inb => n142, outb => n1895);
   U178 : aoi22 port map( a => n143, b => top_data(16), c => n144, d => 
                           load_n_store_lazy_in_2_0_port, outb => n142);
   U179 : inv port map( inb => n145, outb => n1896);
   U180 : aoi22 port map( a => n143, b => top_data(17), c => n144, d => 
                           load_n_store_lazy_in_2_1_port, outb => n145);
   U181 : inv port map( inb => n146, outb => n1897);
   U182 : aoi22 port map( a => n143, b => top_data(18), c => n144, d => 
                           load_n_store_lazy_in_2_2_port, outb => n146);
   U183 : inv port map( inb => n147, outb => n1898);
   U184 : aoi22 port map( a => n143, b => top_data(19), c => n144, d => 
                           load_n_store_lazy_in_2_3_port, outb => n147);
   U185 : inv port map( inb => n148, outb => n1899);
   U186 : aoi22 port map( a => n143, b => top_data(20), c => n144, d => 
                           load_n_store_lazy_in_2_4_port, outb => n148);
   U187 : inv port map( inb => n149, outb => n1900);
   U188 : aoi22 port map( a => n143, b => top_data(21), c => n144, d => 
                           load_n_store_lazy_in_2_5_port, outb => n149);
   U189 : inv port map( inb => n150, outb => n1901);
   U190 : aoi22 port map( a => n143, b => top_data(22), c => n144, d => 
                           load_n_store_lazy_in_2_6_port, outb => n150);
   U191 : inv port map( inb => n151, outb => n1902);
   U192 : aoi22 port map( a => n143, b => top_data(23), c => n144, d => 
                           load_n_store_lazy_in_2_7_port, outb => n151);
   U193 : inv port map( inb => n152, outb => n1903);
   U194 : aoi22 port map( a => n143, b => top_data(8), c => n144, d => 
                           load_n_store_lazy_in_1_0_port, outb => n152);
   U195 : inv port map( inb => n153, outb => n1904);
   U196 : aoi22 port map( a => n143, b => top_data(9), c => n144, d => 
                           load_n_store_lazy_in_1_1_port, outb => n153);
   U197 : inv port map( inb => n154, outb => n1905);
   U198 : aoi22 port map( a => n143, b => top_data(10), c => n144, d => 
                           load_n_store_lazy_in_1_2_port, outb => n154);
   U199 : inv port map( inb => n155, outb => n1906);
   U200 : aoi22 port map( a => n143, b => top_data(11), c => n144, d => 
                           load_n_store_lazy_in_1_3_port, outb => n155);
   U201 : inv port map( inb => n156, outb => n1907);
   U202 : aoi22 port map( a => n143, b => top_data(12), c => n144, d => 
                           load_n_store_lazy_in_1_4_port, outb => n156);
   U203 : inv port map( inb => n157, outb => n1908);
   U204 : aoi22 port map( a => n143, b => top_data(13), c => n144, d => 
                           load_n_store_lazy_in_1_5_port, outb => n157);
   U205 : inv port map( inb => n158, outb => n1909);
   U206 : aoi22 port map( a => n143, b => top_data(14), c => n144, d => 
                           load_n_store_lazy_in_1_6_port, outb => n158);
   U207 : inv port map( inb => n159, outb => n1910);
   U208 : aoi22 port map( a => n143, b => top_data(15), c => n144, d => 
                           load_n_store_lazy_in_1_7_port, outb => n159);
   U209 : inv port map( inb => n160, outb => n1911);
   U210 : aoi22 port map( a => n143, b => top_data(0), c => n144, d => 
                           load_n_store_lazy_in_0_0_port, outb => n160);
   U211 : inv port map( inb => n161, outb => n1912);
   U212 : aoi22 port map( a => n143, b => top_data(1), c => n144, d => 
                           load_n_store_lazy_in_0_1_port, outb => n161);
   U213 : inv port map( inb => n162, outb => n1913);
   U214 : aoi22 port map( a => n143, b => top_data(2), c => n144, d => 
                           load_n_store_lazy_in_0_2_port, outb => n162);
   U215 : inv port map( inb => n163, outb => n1914);
   U216 : aoi22 port map( a => n143, b => top_data(3), c => n144, d => 
                           load_n_store_lazy_in_0_3_port, outb => n163);
   U217 : inv port map( inb => n164, outb => n1915);
   U218 : aoi22 port map( a => n143, b => top_data(4), c => n144, d => 
                           load_n_store_lazy_in_0_4_port, outb => n164);
   U219 : inv port map( inb => n165, outb => n1916);
   U220 : aoi22 port map( a => n143, b => top_data(5), c => n144, d => 
                           load_n_store_lazy_in_0_5_port, outb => n165);
   U221 : inv port map( inb => n166, outb => n1917);
   U222 : aoi22 port map( a => n143, b => top_data(6), c => n144, d => 
                           load_n_store_lazy_in_0_6_port, outb => n166);
   U223 : inv port map( inb => n167, outb => n1918);
   U224 : aoi22 port map( a => n143, b => top_data(7), c => n144, d => 
                           load_n_store_lazy_in_0_7_port, outb => n167);
   U225 : inv port map( inb => n143, outb => n144);
   U226 : nor3 port map( a => n168, b => n169, c => n170, outb => n143);
   U227 : aoi12 port map( b => n171, c => n172, a => n173, outb => n1919);
   U228 : nand2 port map( a => n174, b => n175, outb => n172);
   U229 : oai22 port map( a => n176, b => n177, c => 
                           load_n_store_mem_timer_0_port, d => n178, outb => 
                           n1920);
   U230 : oai12 port map( b => n179, c => n180, a => n181, outb => n1921);
   U231 : nand3 port map( a => n174, b => load_n_store_mem_timer_0_port, c => 
                           n180, outb => n181);
   U232 : oai12 port map( b => n182, c => n183, a => n184, outb => n1922);
   U233 : nand4 port map( a => load_n_store_mem_timer_1_port, b => 
                           load_n_store_mem_timer_0_port, c => n174, d => n183,
                           outb => n184);
   U234 : aoi12 port map( b => n174, c => n180, a => n185, outb => n182);
   U235 : inv port map( inb => n179, outb => n185);
   U236 : aoi12 port map( b => n177, c => n174, a => n186, outb => n179);
   U237 : oai12 port map( b => n187, c => n188, a => n189, outb => n1923);
   U238 : nand3 port map( a => n174, b => n190, c => n188, outb => n189);
   U239 : oai12 port map( b => n191, c => n192, a => n193, outb => n1924);
   U240 : nand4 port map( a => load_n_store_mem_timer_3_port, b => n190, c => 
                           n174, d => n192, outb => n193);
   U241 : aoi12 port map( b => n174, c => n188, a => n194, outb => n191);
   U242 : inv port map( inb => n187, outb => n194);
   U243 : aoi12 port map( b => n195, c => n174, a => n186, outb => n187);
   U244 : oai12 port map( b => n196, c => n197, a => n198, outb => n1925);
   U245 : nand3 port map( a => n174, b => n199, c => n197, outb => n198);
   U246 : oai12 port map( b => n200, c => n201, a => n202, outb => n1926);
   U247 : nand4 port map( a => load_n_store_mem_timer_5_port, b => n199, c => 
                           n174, d => n201, outb => n202);
   U248 : aoi12 port map( b => n174, c => n197, a => n203, outb => n200);
   U249 : inv port map( inb => n196, outb => n203);
   U250 : aoi12 port map( b => n204, c => n174, a => n186, outb => n196);
   U251 : oai12 port map( b => n205, c => n206, a => n207, outb => n1927);
   U252 : nand3 port map( a => n174, b => n208, c => n206, outb => n207);
   U253 : oai12 port map( b => n209, c => n210, a => n211, outb => n1928);
   U254 : nand4 port map( a => load_n_store_mem_timer_7_port, b => n208, c => 
                           n174, d => n210, outb => n211);
   U255 : aoi12 port map( b => n174, c => n206, a => n212, outb => n209);
   U256 : inv port map( inb => n205, outb => n212);
   U257 : aoi12 port map( b => n213, c => n174, a => n186, outb => n205);
   U258 : oai12 port map( b => n214, c => n215, a => n216, outb => n1929);
   U259 : nand3 port map( a => n174, b => n217, c => n215, outb => n216);
   U260 : oai12 port map( b => n218, c => n219, a => n220, outb => n1930);
   U261 : nand4 port map( a => load_n_store_mem_timer_9_port, b => n217, c => 
                           n174, d => n219, outb => n220);
   U262 : aoi12 port map( b => n174, c => n215, a => n221, outb => n218);
   U263 : inv port map( inb => n214, outb => n221);
   U264 : aoi12 port map( b => n222, c => n174, a => n186, outb => n214);
   U265 : oai12 port map( b => n223, c => n224, a => n225, outb => n1931);
   U266 : nand3 port map( a => n174, b => n226, c => n224, outb => n225);
   U267 : oai12 port map( b => n227, c => n228, a => n229, outb => n1932);
   U268 : nand4 port map( a => load_n_store_mem_timer_11_port, b => n226, c => 
                           n174, d => n228, outb => n229);
   U269 : aoi12 port map( b => n174, c => n224, a => n230, outb => n227);
   U270 : inv port map( inb => n223, outb => n230);
   U271 : aoi12 port map( b => n231, c => n174, a => n186, outb => n223);
   U272 : oai12 port map( b => n232, c => n233, a => n234, outb => n1933);
   U273 : nand3 port map( a => n174, b => n235, c => n233, outb => n234);
   U274 : oai12 port map( b => n236, c => n237, a => n238, outb => n1934);
   U275 : nand4 port map( a => load_n_store_mem_timer_13_port, b => n235, c => 
                           n174, d => n237, outb => n238);
   U276 : aoi12 port map( b => n174, c => n233, a => n239, outb => n236);
   U277 : inv port map( inb => n232, outb => n239);
   U278 : aoi12 port map( b => n240, c => n174, a => n186, outb => n232);
   U279 : oai12 port map( b => n241, c => n242, a => n243, outb => n1935);
   U280 : nand3 port map( a => n174, b => n244, c => n242, outb => n243);
   U281 : oai12 port map( b => n245, c => n246, a => n247, outb => n1936);
   U282 : nand4 port map( a => load_n_store_mem_timer_15_port, b => n244, c => 
                           n174, d => n246, outb => n247);
   U283 : aoi12 port map( b => n174, c => n242, a => n248, outb => n245);
   U284 : inv port map( inb => n241, outb => n248);
   U285 : aoi12 port map( b => n249, c => n174, a => n186, outb => n241);
   U286 : oai12 port map( b => n250, c => n251, a => n252, outb => n1937);
   U287 : nand3 port map( a => n174, b => n253, c => n251, outb => n252);
   U288 : oai12 port map( b => n254, c => n255, a => n256, outb => n1938);
   U289 : nand4 port map( a => load_n_store_mem_timer_17_port, b => n253, c => 
                           n174, d => n255, outb => n256);
   U290 : aoi12 port map( b => n174, c => n251, a => n257, outb => n254);
   U291 : inv port map( inb => n250, outb => n257);
   U292 : aoi12 port map( b => n258, c => n174, a => n186, outb => n250);
   U293 : oai12 port map( b => n259, c => n260, a => n261, outb => n1939);
   U294 : nand3 port map( a => n174, b => n262, c => n260, outb => n261);
   U295 : oai12 port map( b => n263, c => n264, a => n265, outb => n1940);
   U296 : nand4 port map( a => load_n_store_mem_timer_19_port, b => n262, c => 
                           n174, d => n264, outb => n265);
   U297 : aoi12 port map( b => n174, c => n260, a => n266, outb => n263);
   U298 : inv port map( inb => n259, outb => n266);
   U299 : aoi12 port map( b => n267, c => n174, a => n186, outb => n259);
   U300 : oai12 port map( b => n268, c => n269, a => n270, outb => n1941);
   U301 : nand3 port map( a => n174, b => n271, c => n269, outb => n270);
   U302 : oai12 port map( b => n272, c => n273, a => n274, outb => n1942);
   U303 : nand4 port map( a => load_n_store_mem_timer_21_port, b => n271, c => 
                           n174, d => n273, outb => n274);
   U304 : aoi12 port map( b => n174, c => n269, a => n275, outb => n272);
   U305 : inv port map( inb => n268, outb => n275);
   U306 : aoi12 port map( b => n276, c => n174, a => n186, outb => n268);
   U307 : oai12 port map( b => n277, c => n278, a => n279, outb => n1943);
   U308 : nand3 port map( a => n174, b => n280, c => n278, outb => n279);
   U309 : oai12 port map( b => n281, c => n282, a => n283, outb => n1944);
   U310 : nand4 port map( a => load_n_store_mem_timer_23_port, b => n280, c => 
                           n174, d => n282, outb => n283);
   U311 : aoi12 port map( b => n174, c => n278, a => n284, outb => n281);
   U312 : inv port map( inb => n277, outb => n284);
   U313 : aoi12 port map( b => n285, c => n174, a => n186, outb => n277);
   U314 : oai12 port map( b => n286, c => n287, a => n288, outb => n1945);
   U315 : nand3 port map( a => n174, b => n289, c => n287, outb => n288);
   U316 : inv port map( inb => n290, outb => n286);
   U317 : oai12 port map( b => n291, c => n292, a => n293, outb => n1946);
   U318 : nand4 port map( a => load_n_store_mem_timer_25_port, b => n289, c => 
                           n174, d => n292, outb => n293);
   U319 : inv port map( inb => load_n_store_mem_timer_26_port, outb => n292);
   U320 : aoi12 port map( b => n174, c => n287, a => n290, outb => n291);
   U321 : oai12 port map( b => n289, c => n178, a => n176, outb => n290);
   U322 : inv port map( inb => load_n_store_mem_timer_25_port, outb => n287);
   U323 : oai12 port map( b => n294, c => n295, a => n296, outb => n1947);
   U324 : nand3 port map( a => n174, b => n297, c => n295, outb => n296);
   U325 : oai12 port map( b => n298, c => n299, a => n300, outb => n1948);
   U326 : nand4 port map( a => load_n_store_mem_timer_27_port, b => n297, c => 
                           n174, d => n299, outb => n300);
   U327 : inv port map( inb => n301, outb => n297);
   U328 : aoi12 port map( b => n174, c => n295, a => n302, outb => n298);
   U329 : inv port map( inb => n294, outb => n302);
   U330 : aoi12 port map( b => n301, c => n174, a => n186, outb => n294);
   U331 : oai12 port map( b => n303, c => n304, a => n305, outb => n1949);
   U332 : nand3 port map( a => n306, b => n174, c => n304, outb => n305);
   U333 : inv port map( inb => n307, outb => n303);
   U334 : oai12 port map( b => n171, c => n175, a => n308, outb => n1950);
   U335 : nand4 port map( a => n306, b => n174, c => 
                           load_n_store_mem_timer_29_port, d => n175, outb => 
                           n308);
   U336 : aoi12 port map( b => n304, c => n174, a => n307, outb => n171);
   U337 : oai12 port map( b => n306, c => n178, a => n176, outb => n307);
   U338 : inv port map( inb => n186, outb => n176);
   U339 : inv port map( inb => n174, outb => n178);
   U340 : nor3 port map( a => n295, b => n301, c => n299, outb => n306);
   U341 : nand3 port map( a => load_n_store_mem_timer_25_port, b => n289, c => 
                           load_n_store_mem_timer_26_port, outb => n301);
   U342 : nor3 port map( a => n278, b => n285, c => n282, outb => n289);
   U343 : inv port map( inb => load_n_store_mem_timer_24_port, outb => n282);
   U344 : inv port map( inb => n280, outb => n285);
   U345 : nor3 port map( a => n269, b => n276, c => n273, outb => n280);
   U346 : inv port map( inb => load_n_store_mem_timer_22_port, outb => n273);
   U347 : inv port map( inb => n271, outb => n276);
   U348 : nor3 port map( a => n260, b => n267, c => n264, outb => n271);
   U349 : inv port map( inb => n262, outb => n267);
   U350 : nor3 port map( a => n251, b => n258, c => n255, outb => n262);
   U351 : inv port map( inb => load_n_store_mem_timer_18_port, outb => n255);
   U352 : inv port map( inb => n253, outb => n258);
   U353 : nor3 port map( a => n242, b => n249, c => n246, outb => n253);
   U354 : inv port map( inb => load_n_store_mem_timer_16_port, outb => n246);
   U355 : inv port map( inb => n244, outb => n249);
   U356 : nor3 port map( a => n233, b => n240, c => n237, outb => n244);
   U357 : inv port map( inb => n235, outb => n240);
   U358 : nor3 port map( a => n224, b => n231, c => n228, outb => n235);
   U359 : inv port map( inb => n226, outb => n231);
   U360 : nor3 port map( a => n219, b => n222, c => n215, outb => n226);
   U361 : inv port map( inb => n217, outb => n222);
   U362 : nor3 port map( a => n206, b => n213, c => n210, outb => n217);
   U363 : inv port map( inb => n208, outb => n213);
   U364 : nor3 port map( a => n197, b => n204, c => n201, outb => n208);
   U365 : inv port map( inb => n199, outb => n204);
   U366 : nor3 port map( a => n188, b => n195, c => n192, outb => n199);
   U367 : inv port map( inb => load_n_store_mem_timer_17_port, outb => n251);
   U368 : inv port map( inb => load_n_store_mem_timer_21_port, outb => n269);
   U369 : inv port map( inb => load_n_store_mem_timer_23_port, outb => n278);
   U370 : inv port map( inb => load_n_store_mem_timer_27_port, outb => n295);
   U371 : nor2 port map( a => n309, b => n186, outb => n174);
   U372 : oai12 port map( b => n310, c => n311, a => reset_port, outb => n186);
   U373 : inv port map( inb => n312, outb => n1951);
   U374 : aoi22 port map( a => n313, b => load_n_store_lazy_out_2_0_port, c => 
                           n314, d => mem_out_r0_0_port, outb => n312);
   U375 : inv port map( inb => n315, outb => n1952);
   U376 : aoi22 port map( a => n313, b => load_n_store_lazy_out_2_1_port, c => 
                           n314, d => mem_out_r0_1_port, outb => n315);
   U377 : inv port map( inb => n316, outb => n1953);
   U378 : aoi22 port map( a => n313, b => load_n_store_lazy_out_2_2_port, c => 
                           n314, d => mem_out_r0_2_port, outb => n316);
   U379 : inv port map( inb => n317, outb => n1954);
   U380 : aoi22 port map( a => n313, b => load_n_store_lazy_out_2_3_port, c => 
                           n314, d => mem_out_r0_3_port, outb => n317);
   U381 : inv port map( inb => n318, outb => n1955);
   U382 : aoi22 port map( a => n313, b => load_n_store_lazy_out_2_4_port, c => 
                           n314, d => mem_out_r0_4_port, outb => n318);
   U383 : inv port map( inb => n319, outb => n1956);
   U384 : aoi22 port map( a => n313, b => load_n_store_lazy_out_2_5_port, c => 
                           n314, d => mem_out_r0_5_port, outb => n319);
   U385 : inv port map( inb => n320, outb => n1957);
   U386 : aoi22 port map( a => n313, b => load_n_store_lazy_out_2_6_port, c => 
                           n314, d => mem_out_r0_6_port, outb => n320);
   U387 : inv port map( inb => n321, outb => n1958);
   U388 : aoi22 port map( a => n313, b => load_n_store_lazy_out_2_7_port, c => 
                           n314, d => mem_out_r0_7_port, outb => n321);
   U389 : inv port map( inb => n322, outb => n1959);
   U390 : aoi22 port map( a => n313, b => load_n_store_lazy_out_1_0_port, c => 
                           n314, d => mem_out_g0_0_port, outb => n322);
   U391 : inv port map( inb => n323, outb => n1960);
   U392 : aoi22 port map( a => n313, b => load_n_store_lazy_out_1_1_port, c => 
                           n314, d => mem_out_g0_1_port, outb => n323);
   U393 : inv port map( inb => n324, outb => n1961);
   U394 : aoi22 port map( a => n313, b => load_n_store_lazy_out_1_2_port, c => 
                           n314, d => mem_out_g0_2_port, outb => n324);
   U395 : inv port map( inb => n325, outb => n1962);
   U396 : aoi22 port map( a => n313, b => load_n_store_lazy_out_1_3_port, c => 
                           n314, d => mem_out_g0_3_port, outb => n325);
   U397 : inv port map( inb => n326, outb => n1963);
   U398 : aoi22 port map( a => n313, b => load_n_store_lazy_out_1_4_port, c => 
                           n314, d => mem_out_g0_4_port, outb => n326);
   U399 : inv port map( inb => n327, outb => n1964);
   U400 : aoi22 port map( a => n313, b => load_n_store_lazy_out_1_5_port, c => 
                           n314, d => mem_out_g0_5_port, outb => n327);
   U401 : inv port map( inb => n328, outb => n1965);
   U402 : aoi22 port map( a => n313, b => load_n_store_lazy_out_1_6_port, c => 
                           n314, d => mem_out_g0_6_port, outb => n328);
   U403 : inv port map( inb => n329, outb => n1966);
   U404 : aoi22 port map( a => n313, b => load_n_store_lazy_out_1_7_port, c => 
                           n314, d => mem_out_g0_7_port, outb => n329);
   U405 : inv port map( inb => n330, outb => n1967);
   U406 : aoi22 port map( a => n313, b => load_n_store_lazy_out_0_0_port, c => 
                           n314, d => mem_out_b0_0_port, outb => n330);
   U407 : inv port map( inb => n331, outb => n1968);
   U408 : aoi22 port map( a => n313, b => load_n_store_lazy_out_0_1_port, c => 
                           n314, d => mem_out_b0_1_port, outb => n331);
   U409 : inv port map( inb => n332, outb => n1969);
   U410 : aoi22 port map( a => n313, b => load_n_store_lazy_out_0_2_port, c => 
                           n314, d => mem_out_b0_2_port, outb => n332);
   U411 : inv port map( inb => n333, outb => n1970);
   U412 : aoi22 port map( a => n313, b => load_n_store_lazy_out_0_3_port, c => 
                           n314, d => mem_out_b0_3_port, outb => n333);
   U413 : inv port map( inb => n334, outb => n1971);
   U414 : aoi22 port map( a => n313, b => load_n_store_lazy_out_0_4_port, c => 
                           n314, d => mem_out_b0_4_port, outb => n334);
   U415 : inv port map( inb => n335, outb => n1972);
   U416 : aoi22 port map( a => n313, b => load_n_store_lazy_out_0_5_port, c => 
                           n314, d => mem_out_b0_5_port, outb => n335);
   U417 : inv port map( inb => n336, outb => n1973);
   U418 : aoi22 port map( a => n313, b => load_n_store_lazy_out_0_6_port, c => 
                           n314, d => mem_out_b0_6_port, outb => n336);
   U419 : inv port map( inb => n337, outb => n1974);
   U420 : aoi22 port map( a => n313, b => load_n_store_lazy_out_0_7_port, c => 
                           n314, d => mem_out_b0_7_port, outb => n337);
   U421 : inv port map( inb => n313, outb => n314);
   U422 : nor3 port map( a => n170, b => top_dv_i, c => n338, outb => n313);
   U423 : oai22 port map( a => n128, b => n339, c => n340, d => n341, outb => 
                           n1975);
   U424 : inv port map( inb => display_out_hub_piso_g0_7_port, outb => n341);
   U425 : inv port map( inb => mem_sipo_g0_7_port, outb => n128);
   U426 : oai22 port map( a => n120, b => n339, c => n340, d => n342, outb => 
                           n1976);
   U427 : inv port map( inb => display_out_hub_piso_r0_7_port, outb => n342);
   U428 : inv port map( inb => mem_sipo_r0_7_port, outb => n120);
   U429 : oai22 port map( a => n71, b => n339, c => n340, d => n343, outb => 
                           n1977);
   U430 : inv port map( inb => display_out_hub_piso_b0_7_port, outb => n343);
   U431 : inv port map( inb => n339, outb => n340);
   U432 : inv port map( inb => mem_sipo_b0_7_port, outb => n71);
   U433 : oai22 port map( a => n344, b => n345, c => n346, d => n13, outb => 
                           n1978);
   U434 : nor3 port map( a => n347, b => n19, c => n49, outb => n345);
   U435 : nor2 port map( a => n58, b => n348, outb => n49);
   U436 : nor2 port map( a => n59, b => n51, outb => n19);
   U437 : nor2 port map( a => n17, b => n14, outb => n51);
   U438 : inv port map( inb => registers_reg_col_inc_0_port, outb => n14);
   U439 : inv port map( inb => registers_reg_col_inc_1_port, outb => n17);
   U440 : inv port map( inb => n50, outb => n59);
   U441 : nor2 port map( a => n348, b => n6, outb => n50);
   U442 : nor3 port map( a => n56, b => n10, c => n348, outb => n347);
   U443 : inv port map( inb => n13, outb => n344);
   U444 : nand3 port map( a => n58, b => n6, c => n349, outb => n13);
   U445 : nand2 port map( a => n9, b => n55, outb => n349);
   U446 : inv port map( inb => n10, outb => n55);
   U447 : nand2 port map( a => registers_mem_to_reg_1_port, b => n346, outb => 
                           n10);
   U448 : inv port map( inb => n57, outb => n9);
   U449 : nand2 port map( a => n8, b => n3, outb => n57);
   U450 : inv port map( inb => registers_s_delay_0_port, outb => n3);
   U451 : inv port map( inb => registers_s_delay_1_port, outb => n8);
   U452 : inv port map( inb => n5, outb => n6);
   U453 : nor2 port map( a => n346, b => registers_mem_to_reg_1_port, outb => 
                           n5);
   U454 : inv port map( inb => registers_mem_to_reg_0_port, outb => n346);
   U455 : inv port map( inb => n350, outb => n58);
   U456 : nor2 port map( a => registers_mem_to_reg_1_port, b => 
                           registers_mem_to_reg_0_port, outb => n350);
   U457 : oai22 port map( a => n351, b => n352, c => n353, d => n354, outb => 
                           n1979);
   U458 : aoi12 port map( b => display_out_disp_timer_30_port, c => n355, a => 
                           n356, outb => n353);
   U459 : oai22 port map( a => n357, b => n358, c => n359, d => n360, outb => 
                           n1980);
   U460 : inv port map( inb => display_out_h_row_10_port, outb => n357);
   U461 : oai22 port map( a => n358, b => n361, c => n360, d => n362, outb => 
                           n1981);
   U462 : inv port map( inb => display_out_h_row_11_port, outb => n361);
   U463 : oai22 port map( a => n358, b => n363, c => n364, d => n360, outb => 
                           n1982);
   U464 : inv port map( inb => display_out_h_row_12_port, outb => n363);
   U465 : oai22 port map( a => n358, b => n365, c => n366, d => n360, outb => 
                           n1983);
   U466 : inv port map( inb => display_out_h_row_13_port, outb => n365);
   U467 : oai22 port map( a => n358, b => n367, c => n368, d => n360, outb => 
                           n1984);
   U468 : inv port map( inb => display_out_h_row_14_port, outb => n367);
   U469 : oai22 port map( a => n358, b => n369, c => n370, d => n360, outb => 
                           n1985);
   U470 : inv port map( inb => display_out_h_row_15_port, outb => n369);
   U471 : oai22 port map( a => n358, b => n371, c => n372, d => n360, outb => 
                           n1986);
   U472 : inv port map( inb => display_out_h_row_16_port, outb => n371);
   U473 : oai22 port map( a => n358, b => n373, c => n374, d => n360, outb => 
                           n1987);
   U474 : inv port map( inb => display_out_h_row_17_port, outb => n373);
   U475 : oai22 port map( a => n358, b => n375, c => n376, d => n360, outb => 
                           n1988);
   U476 : inv port map( inb => display_out_h_row_18_port, outb => n375);
   U477 : oai22 port map( a => n358, b => n377, c => n378, d => n360, outb => 
                           n1989);
   U478 : inv port map( inb => display_out_h_row_19_port, outb => n377);
   U479 : oai22 port map( a => n358, b => n379, c => n380, d => n360, outb => 
                           n1990);
   U480 : inv port map( inb => display_out_h_row_20_port, outb => n379);
   U481 : oai22 port map( a => n358, b => n381, c => n382, d => n360, outb => 
                           n1991);
   U482 : inv port map( inb => display_out_h_row_21_port, outb => n381);
   U483 : oai22 port map( a => n358, b => n383, c => n384, d => n360, outb => 
                           n1992);
   U484 : inv port map( inb => display_out_h_row_22_port, outb => n383);
   U485 : oai22 port map( a => n358, b => n385, c => n386, d => n360, outb => 
                           n1993);
   U486 : inv port map( inb => display_out_h_row_23_port, outb => n385);
   U487 : oai22 port map( a => n358, b => n387, c => n388, d => n360, outb => 
                           n1994);
   U488 : inv port map( inb => display_out_h_row_24_port, outb => n387);
   U489 : oai22 port map( a => n358, b => n389, c => n390, d => n360, outb => 
                           n1995);
   U490 : inv port map( inb => display_out_h_row_25_port, outb => n389);
   U491 : oai22 port map( a => n358, b => n391, c => n360, d => n392, outb => 
                           n1996);
   U492 : inv port map( inb => display_out_h_row_26_port, outb => n391);
   U493 : oai22 port map( a => n358, b => n393, c => n394, d => n360, outb => 
                           n1997);
   U494 : inv port map( inb => display_out_h_row_27_port, outb => n393);
   U495 : oai22 port map( a => n358, b => n395, c => n360, d => n396, outb => 
                           n1998);
   U496 : inv port map( inb => display_out_h_row_28_port, outb => n395);
   U497 : oai22 port map( a => n358, b => n397, c => n398, d => n360, outb => 
                           n1999);
   U498 : inv port map( inb => display_out_h_row_29_port, outb => n397);
   U499 : oai22 port map( a => n358, b => n399, c => n360, d => n400, outb => 
                           n2000);
   U500 : inv port map( inb => display_out_h_row_30_port, outb => n399);
   U501 : oai22 port map( a => n358, b => n401, c => n402, d => n360, outb => 
                           n2001);
   U502 : inv port map( inb => display_out_h_row_31_port, outb => n401);
   U503 : oai22 port map( a => n403, b => n358, c => n360, d => n404, outb => 
                           n2002);
   U504 : inv port map( inb => display_out_h_row_9_port, outb => n403);
   U505 : oai22 port map( a => n405, b => n358, c => n406, d => n360, outb => 
                           n2003);
   U506 : inv port map( inb => display_out_h_row_8_port, outb => n405);
   U507 : oai22 port map( a => n407, b => n358, c => n360, d => n408, outb => 
                           n2004);
   U508 : inv port map( inb => display_out_h_row_7_port, outb => n407);
   U509 : oai22 port map( a => n409, b => n358, c => n360, d => n410, outb => 
                           n2005);
   U510 : inv port map( inb => display_out_h_row_6_port, outb => n409);
   U511 : oai22 port map( a => n411, b => n358, c => n412, d => n360, outb => 
                           n2006);
   U512 : inv port map( inb => display_out_h_row_5_port, outb => n411);
   U513 : oai22 port map( a => n413, b => n358, c => n360, d => n414, outb => 
                           n2007);
   U514 : inv port map( inb => display_out_h_row_4_port, outb => n413);
   U515 : inv port map( inb => n415, outb => n2008);
   U516 : aoi22 port map( a => display_out_h_row_3_port, b => n416, c => n417, 
                           d => n418, outb => n415);
   U517 : oai22 port map( a => n419, b => n358, c => n420, d => n360, outb => 
                           n2009);
   U518 : inv port map( inb => display_out_h_row_2_port, outb => n419);
   U519 : inv port map( inb => n421, outb => n2010);
   U520 : aoi22 port map( a => display_out_h_row_0_port, b => n416, c => n422, 
                           d => n418, outb => n421);
   U521 : oai22 port map( a => n423, b => n358, c => n360, d => n424, outb => 
                           n2011);
   U522 : inv port map( inb => n418, outb => n360);
   U523 : inv port map( inb => display_out_h_row_1_port, outb => n423);
   U524 : inv port map( inb => n425, outb => n2012);
   U525 : aoi12 port map( b => n356, c => display_out_disp_timer_30_port, a => 
                           n426, outb => n425);
   U526 : nor3 port map( a => n427, b => display_out_disp_timer_29_port, c => 
                           display_out_disp_timer_30_port, outb => n426);
   U527 : oai12 port map( b => n352, c => n428, a => n429, outb => n356);
   U528 : oai22 port map( a => n429, b => n428, c => 
                           display_out_disp_timer_29_port, d => n427, outb => 
                           n2013);
   U529 : aoi12 port map( b => n430, c => n355, a => n431, outb => n429);
   U530 : oai12 port map( b => n432, c => n433, a => n427, outb => n2014);
   U531 : nand2 port map( a => n355, b => n434, outb => n427);
   U532 : aoi12 port map( b => display_out_disp_timer_27_port, c => n355, a => 
                           n435, outb => n432);
   U533 : oai12 port map( b => n436, c => n437, a => n438, outb => n2015);
   U534 : nand3 port map( a => n355, b => n439, c => n437, outb => n438);
   U535 : inv port map( inb => n435, outb => n436);
   U536 : oai12 port map( b => n439, c => n352, a => n440, outb => n435);
   U537 : inv port map( inb => n441, outb => n2016);
   U538 : aoi22 port map( a => n439, b => n355, c => n442, d => 
                           display_out_disp_timer_26_port, outb => n441);
   U539 : oai12 port map( b => n443, c => n352, a => n444, outb => n442);
   U540 : oai12 port map( b => n444, c => n443, a => n445, outb => n2017);
   U541 : inv port map( inb => n446, outb => n445);
   U542 : nor3 port map( a => n352, b => n447, c => 
                           display_out_disp_timer_25_port, outb => n446);
   U543 : inv port map( inb => display_out_disp_timer_25_port, outb => n443);
   U544 : aoi12 port map( b => n355, c => display_out_disp_timer_24_port, a => 
                           n448, outb => n444);
   U545 : oai22 port map( a => n449, b => n450, c => n447, d => n352, outb => 
                           n2018);
   U546 : inv port map( inb => n448, outb => n449);
   U547 : oai12 port map( b => n451, c => n352, a => n440, outb => n448);
   U548 : inv port map( inb => n452, outb => n2019);
   U549 : aoi22 port map( a => n451, b => n355, c => n453, d => 
                           display_out_disp_timer_23_port, outb => n452);
   U550 : oai12 port map( b => n454, c => n352, a => n455, outb => n453);
   U551 : oai12 port map( b => n455, c => n454, a => n456, outb => n2020);
   U552 : inv port map( inb => n457, outb => n456);
   U553 : nor3 port map( a => n352, b => n458, c => 
                           display_out_disp_timer_22_port, outb => n457);
   U554 : inv port map( inb => display_out_disp_timer_22_port, outb => n454);
   U555 : aoi12 port map( b => n458, c => n355, a => n431, outb => n455);
   U556 : oai22 port map( a => n458, b => n352, c => n459, d => n460, outb => 
                           n2021);
   U557 : aoi12 port map( b => display_out_disp_timer_20_port, c => n355, a => 
                           n461, outb => n459);
   U558 : oai12 port map( b => n462, c => n463, a => n464, outb => n2022);
   U559 : nand3 port map( a => n355, b => n465, c => n463, outb => n464);
   U560 : inv port map( inb => n461, outb => n462);
   U561 : oai12 port map( b => n465, c => n352, a => n440, outb => n461);
   U562 : inv port map( inb => n466, outb => n2023);
   U563 : aoi22 port map( a => n465, b => n355, c => n467, d => 
                           display_out_disp_timer_19_port, outb => n466);
   U564 : oai12 port map( b => n468, c => n352, a => n469, outb => n467);
   U565 : oai12 port map( b => n469, c => n468, a => n470, outb => n2024);
   U566 : nand3 port map( a => n355, b => n471, c => n468, outb => n470);
   U567 : inv port map( inb => display_out_disp_timer_18_port, outb => n468);
   U568 : aoi12 port map( b => n472, c => n355, a => n431, outb => n469);
   U569 : inv port map( inb => n473, outb => n2025);
   U570 : aoi22 port map( a => n471, b => n355, c => n474, d => 
                           display_out_disp_timer_17_port, outb => n473);
   U571 : oai12 port map( b => n475, c => n352, a => n476, outb => n474);
   U572 : oai12 port map( b => n476, c => n475, a => n477, outb => n2026);
   U573 : nand3 port map( a => n355, b => n478, c => n475, outb => n477);
   U574 : inv port map( inb => n479, outb => n478);
   U575 : aoi12 port map( b => n479, c => n355, a => n431, outb => n476);
   U576 : oai22 port map( a => n479, b => n352, c => n480, d => n481, outb => 
                           n2027);
   U577 : aoi12 port map( b => display_out_disp_timer_14_port, c => n355, a => 
                           n482, outb => n480);
   U578 : oai12 port map( b => n483, c => n484, a => n485, outb => n2028);
   U579 : nand3 port map( a => n355, b => n486, c => n484, outb => n485);
   U580 : inv port map( inb => n482, outb => n483);
   U581 : oai12 port map( b => n486, c => n352, a => n440, outb => n482);
   U582 : nand2 port map( a => n487, b => n488, outb => load_n_store_n303);
   U583 : nand3 port map( a => n310, b => n168, c => reset_port, outb => n487);
   U584 : oai22 port map( a => n489, b => n490, c => n491, d => n488, outb => 
                           load_n_store_n302);
   U585 : nor3 port map( a => n492, b => n493, c => n311, outb => n490);
   U586 : oai12 port map( b => n494, c => n309, a => reset_port, outb => n492);
   U587 : inv port map( inb => n488, outb => n489);
   U588 : nand4 port map( a => reset_port, b => n495, c => n169, d => n494, 
                           outb => n488);
   U589 : inv port map( inb => n310, outb => n494);
   U590 : nand2 port map( a => n493, b => top_dv_i, outb => n495);
   U591 : inv port map( inb => n338, outb => n493);
   U592 : inv port map( inb => n496, outb => load_n_store_n301);
   U593 : aoi22 port map( a => n497, b => top_ack_port, c => n498, d => n499, 
                           outb => n496);
   U594 : inv port map( inb => n498, outb => n497);
   U595 : oai22 port map( a => n170, b => n141, c => n139, d => n500, outb => 
                           n498);
   U596 : nand3 port map( a => n310, b => top_dv_i, c => reset_port, outb => 
                           n139);
   U597 : inv port map( inb => n311, outb => n141);
   U598 : nor2 port map( a => n169, b => top_dv_i, outb => n311);
   U599 : inv port map( inb => n499, outb => n169);
   U600 : nor2 port map( a => load_n_store_simple_mem_sm_0_port, b => 
                           load_n_store_simple_mem_sm_1_port, outb => n499);
   U601 : oai12 port map( b => n501, c => n502, a => n503, outb => 
                           load_n_store_n300);
   U602 : oai12 port map( b => n348, c => n502, a => n503, outb => 
                           load_n_store_n299);
   U603 : nand3 port map( a => n502, b => n168, c => reset_port, outb => n503);
   U604 : inv port map( inb => top_dv_i, outb => n168);
   U605 : nand2 port map( a => n140, b => n338, outb => n502);
   U606 : nand2 port map( a => load_n_store_simple_mem_sm_1_port, b => n491, 
                           outb => n338);
   U607 : aoi12 port map( b => n309, c => n310, a => n170, outb => n140);
   U608 : inv port map( inb => reset_port, outb => n170);
   U609 : nor2 port map( a => n491, b => load_n_store_simple_mem_sm_1_port, 
                           outb => n310);
   U610 : inv port map( inb => load_n_store_simple_mem_sm_0_port, outb => n491)
                           ;
   U611 : nand2 port map( a => top_dv_i, b => n500, outb => n309);
   U612 : nand2 port map( a => n504, b => n173, outb => n500);
   U613 : inv port map( inb => load_n_store_mem_timer_31_port, outb => n173);
   U614 : nand2 port map( a => n505, b => n506, outb => n504);
   U615 : nor3 port map( a => n507, b => n508, c => n509, outb => n506);
   U616 : nand4 port map( a => n175, b => n188, c => n192, d => n197, outb => 
                           n509);
   U617 : inv port map( inb => load_n_store_mem_timer_5_port, outb => n197);
   U618 : inv port map( inb => load_n_store_mem_timer_4_port, outb => n192);
   U619 : inv port map( inb => load_n_store_mem_timer_3_port, outb => n188);
   U620 : inv port map( inb => load_n_store_mem_timer_30_port, outb => n175);
   U621 : nand4 port map( a => n201, b => n206, c => n210, d => n215, outb => 
                           n508);
   U622 : inv port map( inb => load_n_store_mem_timer_9_port, outb => n215);
   U623 : inv port map( inb => load_n_store_mem_timer_8_port, outb => n210);
   U624 : inv port map( inb => load_n_store_mem_timer_7_port, outb => n206);
   U625 : inv port map( inb => load_n_store_mem_timer_6_port, outb => n201);
   U626 : nand4 port map( a => n299, b => n304, c => n510, d => n511, outb => 
                           n507);
   U627 : nor3 port map( a => load_n_store_mem_timer_23_port, b => 
                           load_n_store_mem_timer_25_port, c => 
                           load_n_store_mem_timer_24_port, outb => n511);
   U628 : nor2 port map( a => load_n_store_mem_timer_27_port, b => 
                           load_n_store_mem_timer_26_port, outb => n510);
   U629 : inv port map( inb => load_n_store_mem_timer_29_port, outb => n304);
   U630 : inv port map( inb => load_n_store_mem_timer_28_port, outb => n299);
   U631 : nor3 port map( a => n512, b => n513, c => n514, outb => n505);
   U632 : nand3 port map( a => n219, b => n224, c => n195, outb => n514);
   U633 : inv port map( inb => n190, outb => n195);
   U634 : nor3 port map( a => n180, b => n177, c => n183, outb => n190);
   U635 : inv port map( inb => load_n_store_mem_timer_2_port, outb => n183);
   U636 : inv port map( inb => load_n_store_mem_timer_0_port, outb => n177);
   U637 : inv port map( inb => load_n_store_mem_timer_1_port, outb => n180);
   U638 : inv port map( inb => load_n_store_mem_timer_11_port, outb => n224);
   U639 : inv port map( inb => load_n_store_mem_timer_10_port, outb => n219);
   U640 : nand4 port map( a => n228, b => n233, c => n237, d => n242, outb => 
                           n513);
   U641 : inv port map( inb => load_n_store_mem_timer_15_port, outb => n242);
   U642 : inv port map( inb => load_n_store_mem_timer_14_port, outb => n237);
   U643 : inv port map( inb => load_n_store_mem_timer_13_port, outb => n233);
   U644 : inv port map( inb => load_n_store_mem_timer_12_port, outb => n228);
   U645 : nand4 port map( a => n260, b => n264, c => n515, d => n516, outb => 
                           n512);
   U646 : nor3 port map( a => load_n_store_mem_timer_16_port, b => 
                           load_n_store_mem_timer_18_port, c => 
                           load_n_store_mem_timer_17_port, outb => n516);
   U647 : nor2 port map( a => load_n_store_mem_timer_22_port, b => 
                           load_n_store_mem_timer_21_port, outb => n515);
   U648 : inv port map( inb => load_n_store_mem_timer_20_port, outb => n264);
   U649 : inv port map( inb => load_n_store_mem_timer_19_port, outb => n260);
   U650 : inv port map( inb => mem_reg_f, outb => n348);
   U651 : nand3 port map( a => n517, b => n518, c => n519, outb => n2304);
   U652 : nand2 port map( a => load_n_store_lazy_in_2_3_port, b => 
                           load_n_store_we_i, outb => n519);
   U653 : nand4 port map( a => n520, b => n521, c => n522, d => n523, outb => 
                           n518);
   U654 : nor3 port map( a => n524, b => n525, c => n526, outb => n523);
   U655 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_5_3_port, b
                           => n527, c => 
                           load_n_store_RGB_Array_2_block_ram_r_3_3_port, d => 
                           n528, outb => n526);
   U656 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_7_3_port, b 
                           => n529, outb => n525);
   U657 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_1_3_port, b
                           => n530, c => 
                           load_n_store_RGB_Array_2_block_ram_r_0_3_port, d => 
                           n531, outb => n524);
   U658 : aoi22 port map( a => n532, b => n533, c => n534, d => n535, outb => 
                           n522);
   U659 : nand2 port map( a => n536, b => n537, outb => n521);
   U660 : nand4 port map( a => n538, b => n539, c => n540, d => n541, outb => 
                           n517);
   U661 : nor3 port map( a => n542, b => n543, c => n544, outb => n541);
   U662 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_13_3_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_2_block_ram_r_11_3_port, d =>
                           n528, outb => n544);
   U663 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_15_3_port, b
                           => n529, outb => n543);
   U664 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_9_3_port, b
                           => n530, c => 
                           load_n_store_RGB_Array_2_block_ram_r_8_3_port, d => 
                           n531, outb => n542);
   U665 : aoi22 port map( a => n532, b => n545, c => n534, d => n546, outb => 
                           n540);
   U666 : nand2 port map( a => n536, b => n547, outb => n539);
   U667 : inv port map( inb => n548, outb => n2572);
   U668 : aoi22 port map( a => load_n_store_lazy_in_2_7_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_2_block_ram_r_15_7_port, outb
                           => n548);
   U669 : inv port map( inb => n551, outb => n2571);
   U670 : aoi22 port map( a => load_n_store_lazy_in_2_6_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_2_block_ram_r_15_6_port, outb
                           => n551);
   U671 : inv port map( inb => n552, outb => n2570);
   U672 : aoi22 port map( a => load_n_store_lazy_in_2_5_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_2_block_ram_r_15_5_port, outb
                           => n552);
   U673 : inv port map( inb => n553, outb => n2569);
   U674 : aoi22 port map( a => load_n_store_lazy_in_2_4_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_2_block_ram_r_15_4_port, outb
                           => n553);
   U675 : inv port map( inb => n554, outb => n2568);
   U676 : aoi22 port map( a => load_n_store_lazy_in_2_3_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_2_block_ram_r_15_3_port, outb
                           => n554);
   U677 : inv port map( inb => n555, outb => n2567);
   U678 : aoi22 port map( a => load_n_store_lazy_in_2_2_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_2_block_ram_r_15_2_port, outb
                           => n555);
   U679 : inv port map( inb => n556, outb => n2566);
   U680 : aoi22 port map( a => load_n_store_lazy_in_2_1_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_2_block_ram_r_15_1_port, outb
                           => n556);
   U681 : inv port map( inb => n557, outb => n2565);
   U682 : aoi22 port map( a => load_n_store_lazy_in_2_0_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_2_block_ram_r_15_0_port, outb
                           => n557);
   U683 : oai22 port map( a => n558, b => n559, c => n560, d => n561, outb => 
                           n2564);
   U684 : oai22 port map( a => n562, b => n559, c => n560, d => n563, outb => 
                           n2563);
   U685 : oai22 port map( a => n564, b => n559, c => n560, d => n565, outb => 
                           n2562);
   U686 : nand3 port map( a => n566, b => n567, c => n568, outb => n2303);
   U687 : nand2 port map( a => load_n_store_lazy_in_2_2_port, b => 
                           load_n_store_we_i, outb => n568);
   U688 : nand4 port map( a => n520, b => n569, c => n570, d => n571, outb => 
                           n567);
   U689 : nor3 port map( a => n572, b => n573, c => n574, outb => n571);
   U690 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_5_2_port, b
                           => n527, c => 
                           load_n_store_RGB_Array_2_block_ram_r_3_2_port, d => 
                           n528, outb => n574);
   U691 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_7_2_port, b 
                           => n529, outb => n573);
   U692 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_1_2_port, b
                           => n530, c => 
                           load_n_store_RGB_Array_2_block_ram_r_0_2_port, d => 
                           n531, outb => n572);
   U693 : aoi22 port map( a => n532, b => n575, c => n534, d => n576, outb => 
                           n570);
   U694 : nand2 port map( a => n536, b => n577, outb => n569);
   U695 : nand4 port map( a => n538, b => n578, c => n579, d => n580, outb => 
                           n566);
   U696 : nor3 port map( a => n581, b => n582, c => n583, outb => n580);
   U697 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_13_2_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_2_block_ram_r_11_2_port, d =>
                           n528, outb => n583);
   U698 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_15_2_port, b
                           => n529, outb => n582);
   U699 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_9_2_port, b
                           => n530, c => 
                           load_n_store_RGB_Array_2_block_ram_r_8_2_port, d => 
                           n531, outb => n581);
   U700 : aoi22 port map( a => n532, b => n584, c => n534, d => n585, outb => 
                           n579);
   U701 : nand2 port map( a => n536, b => n586, outb => n578);
   U702 : oai22 port map( a => n587, b => n559, c => n560, d => n588, outb => 
                           n2561);
   U703 : oai22 port map( a => n589, b => n559, c => n560, d => n547, outb => 
                           n2560);
   U704 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_14_3_port, 
                           outb => n547);
   U705 : oai22 port map( a => n590, b => n559, c => n560, d => n586, outb => 
                           n2559);
   U706 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_14_2_port, 
                           outb => n586);
   U707 : oai22 port map( a => n591, b => n559, c => n560, d => n592, outb => 
                           n2558);
   U708 : oai22 port map( a => n593, b => n559, c => n560, d => n594, outb => 
                           n2557);
   U709 : inv port map( inb => n595, outb => n2556);
   U710 : aoi22 port map( a => load_n_store_lazy_in_2_7_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_2_block_ram_r_13_7_port, outb
                           => n595);
   U711 : inv port map( inb => n598, outb => n2555);
   U712 : aoi22 port map( a => load_n_store_lazy_in_2_6_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_2_block_ram_r_13_6_port, outb
                           => n598);
   U713 : inv port map( inb => n599, outb => n2554);
   U714 : aoi22 port map( a => load_n_store_lazy_in_2_5_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_2_block_ram_r_13_5_port, outb
                           => n599);
   U715 : inv port map( inb => n600, outb => n2553);
   U716 : aoi22 port map( a => load_n_store_lazy_in_2_4_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_2_block_ram_r_13_4_port, outb
                           => n600);
   U717 : inv port map( inb => n601, outb => n2552);
   U718 : aoi22 port map( a => load_n_store_lazy_in_2_3_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_2_block_ram_r_13_3_port, outb
                           => n601);
   U719 : inv port map( inb => n602, outb => n2551);
   U720 : aoi22 port map( a => load_n_store_lazy_in_2_2_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_2_block_ram_r_13_2_port, outb
                           => n602);
   U721 : inv port map( inb => n603, outb => n2550);
   U722 : aoi22 port map( a => load_n_store_lazy_in_2_1_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_2_block_ram_r_13_1_port, outb
                           => n603);
   U723 : inv port map( inb => n604, outb => n2549);
   U724 : aoi22 port map( a => load_n_store_lazy_in_2_0_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_2_block_ram_r_13_0_port, outb
                           => n604);
   U725 : oai22 port map( a => n558, b => n605, c => n606, d => n607, outb => 
                           n2548);
   U726 : oai22 port map( a => n562, b => n605, c => n606, d => n608, outb => 
                           n2547);
   U727 : oai22 port map( a => n564, b => n605, c => n606, d => n609, outb => 
                           n2546);
   U728 : oai22 port map( a => n587, b => n605, c => n606, d => n610, outb => 
                           n2545);
   U729 : oai22 port map( a => n589, b => n605, c => n606, d => n545, outb => 
                           n2544);
   U730 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_12_3_port, 
                           outb => n545);
   U731 : oai22 port map( a => n590, b => n605, c => n606, d => n584, outb => 
                           n2543);
   U732 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_12_2_port, 
                           outb => n584);
   U733 : oai22 port map( a => n591, b => n605, c => n606, d => n611, outb => 
                           n2542);
   U734 : oai22 port map( a => n593, b => n605, c => n606, d => n612, outb => 
                           n2541);
   U735 : inv port map( inb => n613, outb => n2540);
   U736 : aoi22 port map( a => load_n_store_lazy_in_2_7_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_2_block_ram_r_11_7_port, outb
                           => n613);
   U737 : inv port map( inb => n616, outb => n2539);
   U738 : aoi22 port map( a => load_n_store_lazy_in_2_6_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_2_block_ram_r_11_6_port, outb
                           => n616);
   U739 : inv port map( inb => n617, outb => n2538);
   U740 : aoi22 port map( a => load_n_store_lazy_in_2_5_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_2_block_ram_r_11_5_port, outb
                           => n617);
   U741 : inv port map( inb => n618, outb => n2537);
   U742 : aoi22 port map( a => load_n_store_lazy_in_2_4_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_2_block_ram_r_11_4_port, outb
                           => n618);
   U743 : inv port map( inb => n619, outb => n2536);
   U744 : aoi22 port map( a => load_n_store_lazy_in_2_3_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_2_block_ram_r_11_3_port, outb
                           => n619);
   U745 : inv port map( inb => n620, outb => n2535);
   U746 : aoi22 port map( a => load_n_store_lazy_in_2_2_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_2_block_ram_r_11_2_port, outb
                           => n620);
   U747 : inv port map( inb => n621, outb => n2534);
   U748 : aoi22 port map( a => load_n_store_lazy_in_2_1_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_2_block_ram_r_11_1_port, outb
                           => n621);
   U749 : inv port map( inb => n622, outb => n2533);
   U750 : aoi22 port map( a => load_n_store_lazy_in_2_0_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_2_block_ram_r_11_0_port, outb
                           => n622);
   U751 : oai22 port map( a => n558, b => n623, c => n624, d => n625, outb => 
                           n2532);
   U752 : oai22 port map( a => n562, b => n623, c => n624, d => n626, outb => 
                           n2531);
   U753 : oai22 port map( a => n564, b => n623, c => n624, d => n627, outb => 
                           n2530);
   U754 : oai22 port map( a => n587, b => n623, c => n624, d => n628, outb => 
                           n2529);
   U755 : oai22 port map( a => n589, b => n623, c => n624, d => n546, outb => 
                           n2528);
   U756 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_10_3_port, 
                           outb => n546);
   U757 : oai22 port map( a => n590, b => n623, c => n624, d => n585, outb => 
                           n2527);
   U758 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_10_2_port, 
                           outb => n585);
   U759 : oai22 port map( a => n591, b => n623, c => n624, d => n629, outb => 
                           n2526);
   U760 : oai22 port map( a => n593, b => n623, c => n624, d => n630, outb => 
                           n2525);
   U761 : inv port map( inb => n631, outb => n2524);
   U762 : aoi22 port map( a => load_n_store_lazy_in_2_7_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_2_block_ram_r_9_7_port, outb 
                           => n631);
   U763 : inv port map( inb => n634, outb => n2523);
   U764 : aoi22 port map( a => load_n_store_lazy_in_2_6_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_2_block_ram_r_9_6_port, outb 
                           => n634);
   U765 : inv port map( inb => n635, outb => n2522);
   U766 : aoi22 port map( a => load_n_store_lazy_in_2_5_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_2_block_ram_r_9_5_port, outb 
                           => n635);
   U767 : inv port map( inb => n636, outb => n2521);
   U768 : aoi22 port map( a => load_n_store_lazy_in_2_4_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_2_block_ram_r_9_4_port, outb 
                           => n636);
   U769 : inv port map( inb => n637, outb => n2520);
   U770 : aoi22 port map( a => load_n_store_lazy_in_2_3_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_2_block_ram_r_9_3_port, outb 
                           => n637);
   U771 : inv port map( inb => n638, outb => n2519);
   U772 : aoi22 port map( a => load_n_store_lazy_in_2_2_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_2_block_ram_r_9_2_port, outb 
                           => n638);
   U773 : inv port map( inb => n639, outb => n2518);
   U774 : aoi22 port map( a => load_n_store_lazy_in_2_1_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_2_block_ram_r_9_1_port, outb 
                           => n639);
   U775 : inv port map( inb => n640, outb => n2517);
   U776 : aoi22 port map( a => load_n_store_lazy_in_2_0_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_2_block_ram_r_9_0_port, outb 
                           => n640);
   U777 : inv port map( inb => n641, outb => n2516);
   U778 : aoi22 port map( a => load_n_store_lazy_in_2_7_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_2_block_ram_r_8_7_port, outb 
                           => n641);
   U779 : inv port map( inb => n644, outb => n2515);
   U780 : aoi22 port map( a => load_n_store_lazy_in_2_6_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_2_block_ram_r_8_6_port, outb 
                           => n644);
   U781 : inv port map( inb => n645, outb => n2514);
   U782 : aoi22 port map( a => load_n_store_lazy_in_2_5_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_2_block_ram_r_8_5_port, outb 
                           => n645);
   U783 : inv port map( inb => n646, outb => n2513);
   U784 : aoi22 port map( a => load_n_store_lazy_in_2_4_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_2_block_ram_r_8_4_port, outb 
                           => n646);
   U785 : inv port map( inb => n647, outb => n2512);
   U786 : aoi22 port map( a => load_n_store_lazy_in_2_3_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_2_block_ram_r_8_3_port, outb 
                           => n647);
   U787 : inv port map( inb => n648, outb => n2511);
   U788 : aoi22 port map( a => load_n_store_lazy_in_2_2_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_2_block_ram_r_8_2_port, outb 
                           => n648);
   U789 : inv port map( inb => n649, outb => n2510);
   U790 : aoi22 port map( a => load_n_store_lazy_in_2_1_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_2_block_ram_r_8_1_port, outb 
                           => n649);
   U791 : inv port map( inb => n650, outb => n2509);
   U792 : aoi22 port map( a => load_n_store_lazy_in_2_0_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_2_block_ram_r_8_0_port, outb 
                           => n650);
   U793 : inv port map( inb => n651, outb => n2508);
   U794 : aoi22 port map( a => load_n_store_lazy_in_2_7_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_2_block_ram_r_7_7_port, outb 
                           => n651);
   U795 : inv port map( inb => n654, outb => n2507);
   U796 : aoi22 port map( a => load_n_store_lazy_in_2_6_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_2_block_ram_r_7_6_port, outb 
                           => n654);
   U797 : inv port map( inb => n655, outb => n2506);
   U798 : aoi22 port map( a => load_n_store_lazy_in_2_5_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_2_block_ram_r_7_5_port, outb 
                           => n655);
   U799 : inv port map( inb => n656, outb => n2505);
   U800 : aoi22 port map( a => load_n_store_lazy_in_2_4_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_2_block_ram_r_7_4_port, outb 
                           => n656);
   U801 : inv port map( inb => n657, outb => n2504);
   U802 : aoi22 port map( a => load_n_store_lazy_in_2_3_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_2_block_ram_r_7_3_port, outb 
                           => n657);
   U803 : inv port map( inb => n658, outb => n2503);
   U804 : aoi22 port map( a => load_n_store_lazy_in_2_2_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_2_block_ram_r_7_2_port, outb 
                           => n658);
   U805 : inv port map( inb => n659, outb => n2502);
   U806 : aoi22 port map( a => load_n_store_lazy_in_2_1_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_2_block_ram_r_7_1_port, outb 
                           => n659);
   U807 : inv port map( inb => n660, outb => n2501);
   U808 : aoi22 port map( a => load_n_store_lazy_in_2_0_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_2_block_ram_r_7_0_port, outb 
                           => n660);
   U809 : oai22 port map( a => n558, b => n661, c => n662, d => n663, outb => 
                           n2500);
   U810 : oai22 port map( a => n562, b => n661, c => n662, d => n664, outb => 
                           n2499);
   U811 : oai22 port map( a => n564, b => n661, c => n662, d => n665, outb => 
                           n2498);
   U812 : oai22 port map( a => n587, b => n661, c => n662, d => n666, outb => 
                           n2497);
   U813 : oai22 port map( a => n589, b => n661, c => n662, d => n537, outb => 
                           n2496);
   U814 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_6_3_port, 
                           outb => n537);
   U815 : oai22 port map( a => n590, b => n661, c => n662, d => n577, outb => 
                           n2495);
   U816 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_6_2_port, 
                           outb => n577);
   U817 : oai22 port map( a => n591, b => n661, c => n662, d => n667, outb => 
                           n2494);
   U818 : oai22 port map( a => n593, b => n661, c => n662, d => n668, outb => 
                           n2493);
   U819 : inv port map( inb => n669, outb => n2492);
   U820 : aoi22 port map( a => load_n_store_lazy_in_2_7_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_2_block_ram_r_5_7_port, outb 
                           => n669);
   U821 : inv port map( inb => n672, outb => n2491);
   U822 : aoi22 port map( a => load_n_store_lazy_in_2_6_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_2_block_ram_r_5_6_port, outb 
                           => n672);
   U823 : inv port map( inb => n673, outb => n2490);
   U824 : aoi22 port map( a => load_n_store_lazy_in_2_5_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_2_block_ram_r_5_5_port, outb 
                           => n673);
   U825 : inv port map( inb => n674, outb => n2489);
   U826 : aoi22 port map( a => load_n_store_lazy_in_2_4_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_2_block_ram_r_5_4_port, outb 
                           => n674);
   U827 : inv port map( inb => n675, outb => n2488);
   U828 : aoi22 port map( a => load_n_store_lazy_in_2_3_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_2_block_ram_r_5_3_port, outb 
                           => n675);
   U829 : inv port map( inb => n676, outb => n2487);
   U830 : aoi22 port map( a => load_n_store_lazy_in_2_2_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_2_block_ram_r_5_2_port, outb 
                           => n676);
   U831 : inv port map( inb => n677, outb => n2486);
   U832 : aoi22 port map( a => load_n_store_lazy_in_2_1_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_2_block_ram_r_5_1_port, outb 
                           => n677);
   U833 : inv port map( inb => n678, outb => n2485);
   U834 : aoi22 port map( a => load_n_store_lazy_in_2_0_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_2_block_ram_r_5_0_port, outb 
                           => n678);
   U835 : oai22 port map( a => n558, b => n679, c => n680, d => n681, outb => 
                           n2484);
   U836 : oai22 port map( a => n562, b => n679, c => n680, d => n682, outb => 
                           n2483);
   U837 : oai22 port map( a => n564, b => n679, c => n680, d => n683, outb => 
                           n2482);
   U838 : oai22 port map( a => n587, b => n679, c => n680, d => n684, outb => 
                           n2481);
   U839 : oai22 port map( a => n589, b => n679, c => n680, d => n533, outb => 
                           n2480);
   U840 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_4_3_port, 
                           outb => n533);
   U841 : oai22 port map( a => n590, b => n679, c => n680, d => n575, outb => 
                           n2479);
   U842 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_4_2_port, 
                           outb => n575);
   U843 : oai22 port map( a => n591, b => n679, c => n680, d => n685, outb => 
                           n2478);
   U844 : oai22 port map( a => n593, b => n679, c => n680, d => n686, outb => 
                           n2477);
   U845 : inv port map( inb => n687, outb => n2476);
   U846 : aoi22 port map( a => load_n_store_lazy_in_2_7_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_2_block_ram_r_3_7_port, outb 
                           => n687);
   U847 : inv port map( inb => n690, outb => n2475);
   U848 : aoi22 port map( a => load_n_store_lazy_in_2_6_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_2_block_ram_r_3_6_port, outb 
                           => n690);
   U849 : inv port map( inb => n691, outb => n2474);
   U850 : aoi22 port map( a => load_n_store_lazy_in_2_5_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_2_block_ram_r_3_5_port, outb 
                           => n691);
   U851 : inv port map( inb => n692, outb => n2473);
   U852 : aoi22 port map( a => load_n_store_lazy_in_2_4_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_2_block_ram_r_3_4_port, outb 
                           => n692);
   U853 : inv port map( inb => n693, outb => n2472);
   U854 : aoi22 port map( a => load_n_store_lazy_in_2_3_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_2_block_ram_r_3_3_port, outb 
                           => n693);
   U855 : inv port map( inb => n694, outb => n2471);
   U856 : aoi22 port map( a => load_n_store_lazy_in_2_2_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_2_block_ram_r_3_2_port, outb 
                           => n694);
   U857 : inv port map( inb => n695, outb => n2470);
   U858 : aoi22 port map( a => load_n_store_lazy_in_2_1_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_2_block_ram_r_3_1_port, outb 
                           => n695);
   U859 : inv port map( inb => n696, outb => n2469);
   U860 : aoi22 port map( a => load_n_store_lazy_in_2_0_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_2_block_ram_r_3_0_port, outb 
                           => n696);
   U861 : oai22 port map( a => n558, b => n697, c => n698, d => n699, outb => 
                           n2468);
   U862 : inv port map( inb => load_n_store_lazy_in_2_7_port, outb => n558);
   U863 : oai22 port map( a => n562, b => n697, c => n698, d => n700, outb => 
                           n2467);
   U864 : inv port map( inb => load_n_store_lazy_in_2_6_port, outb => n562);
   U865 : oai22 port map( a => n564, b => n697, c => n698, d => n701, outb => 
                           n2466);
   U866 : inv port map( inb => load_n_store_lazy_in_2_5_port, outb => n564);
   U867 : oai22 port map( a => n587, b => n697, c => n698, d => n702, outb => 
                           n2465);
   U868 : inv port map( inb => load_n_store_lazy_in_2_4_port, outb => n587);
   U869 : oai22 port map( a => n589, b => n697, c => n698, d => n535, outb => 
                           n2464);
   U870 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_2_3_port, 
                           outb => n535);
   U871 : inv port map( inb => load_n_store_lazy_in_2_3_port, outb => n589);
   U872 : oai22 port map( a => n590, b => n697, c => n698, d => n576, outb => 
                           n2463);
   U873 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_2_2_port, 
                           outb => n576);
   U874 : inv port map( inb => load_n_store_lazy_in_2_2_port, outb => n590);
   U875 : oai22 port map( a => n591, b => n697, c => n698, d => n703, outb => 
                           n2462);
   U876 : inv port map( inb => load_n_store_lazy_in_2_1_port, outb => n591);
   U877 : oai22 port map( a => n593, b => n697, c => n698, d => n704, outb => 
                           n2461);
   U878 : inv port map( inb => load_n_store_lazy_in_2_0_port, outb => n593);
   U879 : inv port map( inb => n705, outb => n2460);
   U880 : aoi22 port map( a => load_n_store_lazy_in_2_7_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_2_block_ram_r_1_7_port, outb 
                           => n705);
   U881 : inv port map( inb => n708, outb => n2459);
   U882 : aoi22 port map( a => load_n_store_lazy_in_2_6_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_2_block_ram_r_1_6_port, outb 
                           => n708);
   U883 : inv port map( inb => n709, outb => n2458);
   U884 : aoi22 port map( a => load_n_store_lazy_in_2_5_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_2_block_ram_r_1_5_port, outb 
                           => n709);
   U885 : inv port map( inb => n710, outb => n2457);
   U886 : aoi22 port map( a => load_n_store_lazy_in_2_4_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_2_block_ram_r_1_4_port, outb 
                           => n710);
   U887 : inv port map( inb => n711, outb => n2456);
   U888 : aoi22 port map( a => load_n_store_lazy_in_2_3_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_2_block_ram_r_1_3_port, outb 
                           => n711);
   U889 : inv port map( inb => n712, outb => n2455);
   U890 : aoi22 port map( a => load_n_store_lazy_in_2_2_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_2_block_ram_r_1_2_port, outb 
                           => n712);
   U891 : inv port map( inb => n713, outb => n2454);
   U892 : aoi22 port map( a => load_n_store_lazy_in_2_1_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_2_block_ram_r_1_1_port, outb 
                           => n713);
   U893 : inv port map( inb => n714, outb => n2453);
   U894 : aoi22 port map( a => load_n_store_lazy_in_2_0_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_2_block_ram_r_1_0_port, outb 
                           => n714);
   U895 : inv port map( inb => n715, outb => n2452);
   U896 : aoi22 port map( a => load_n_store_lazy_in_2_7_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_2_block_ram_r_0_7_port, outb 
                           => n715);
   U897 : inv port map( inb => n718, outb => n2451);
   U898 : aoi22 port map( a => load_n_store_lazy_in_2_6_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_2_block_ram_r_0_6_port, outb 
                           => n718);
   U899 : inv port map( inb => n719, outb => n2450);
   U900 : aoi22 port map( a => load_n_store_lazy_in_2_5_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_2_block_ram_r_0_5_port, outb 
                           => n719);
   U901 : inv port map( inb => n720, outb => n2449);
   U902 : aoi22 port map( a => load_n_store_lazy_in_2_4_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_2_block_ram_r_0_4_port, outb 
                           => n720);
   U903 : inv port map( inb => n721, outb => n2448);
   U904 : aoi22 port map( a => load_n_store_lazy_in_2_3_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_2_block_ram_r_0_3_port, outb 
                           => n721);
   U905 : inv port map( inb => n722, outb => n2447);
   U906 : aoi22 port map( a => load_n_store_lazy_in_2_2_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_2_block_ram_r_0_2_port, outb 
                           => n722);
   U907 : inv port map( inb => n723, outb => n2446);
   U908 : aoi22 port map( a => load_n_store_lazy_in_2_1_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_2_block_ram_r_0_1_port, outb 
                           => n723);
   U909 : inv port map( inb => n724, outb => n2445);
   U910 : aoi22 port map( a => load_n_store_lazy_in_2_0_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_2_block_ram_r_0_0_port, outb 
                           => n724);
   U911 : nand3 port map( a => n725, b => n726, c => n727, outb => n2302);
   U912 : nand2 port map( a => load_n_store_lazy_in_2_1_port, b => 
                           load_n_store_we_i, outb => n727);
   U913 : nand4 port map( a => n520, b => n728, c => n729, d => n730, outb => 
                           n726);
   U914 : nor3 port map( a => n731, b => n732, c => n733, outb => n730);
   U915 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_5_1_port, b
                           => n527, c => 
                           load_n_store_RGB_Array_2_block_ram_r_3_1_port, d => 
                           n528, outb => n733);
   U916 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_7_1_port, b 
                           => n529, outb => n732);
   U917 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_1_1_port, b
                           => n530, c => 
                           load_n_store_RGB_Array_2_block_ram_r_0_1_port, d => 
                           n531, outb => n731);
   U918 : aoi22 port map( a => n532, b => n685, c => n534, d => n703, outb => 
                           n729);
   U919 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_2_1_port, 
                           outb => n703);
   U920 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_4_1_port, 
                           outb => n685);
   U921 : nand2 port map( a => n536, b => n667, outb => n728);
   U922 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_6_1_port, 
                           outb => n667);
   U923 : nand4 port map( a => n538, b => n734, c => n735, d => n736, outb => 
                           n725);
   U924 : nor3 port map( a => n737, b => n738, c => n739, outb => n736);
   U925 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_13_1_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_2_block_ram_r_11_1_port, d =>
                           n528, outb => n739);
   U926 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_15_1_port, b
                           => n529, outb => n738);
   U927 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_9_1_port, b
                           => n530, c => 
                           load_n_store_RGB_Array_2_block_ram_r_8_1_port, d => 
                           n531, outb => n737);
   U928 : aoi22 port map( a => n532, b => n611, c => n534, d => n629, outb => 
                           n735);
   U929 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_10_1_port, 
                           outb => n629);
   U930 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_12_1_port, 
                           outb => n611);
   U931 : nand2 port map( a => n536, b => n592, outb => n734);
   U932 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_14_1_port, 
                           outb => n592);
   U933 : nand3 port map( a => n740, b => n741, c => n742, outb => n2301);
   U934 : nand2 port map( a => load_n_store_lazy_in_2_0_port, b => 
                           load_n_store_we_i, outb => n742);
   U935 : nand4 port map( a => n520, b => n743, c => n744, d => n745, outb => 
                           n741);
   U936 : nor3 port map( a => n746, b => n747, c => n748, outb => n745);
   U937 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_5_0_port, b
                           => n527, c => 
                           load_n_store_RGB_Array_2_block_ram_r_3_0_port, d => 
                           n528, outb => n748);
   U938 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_7_0_port, b 
                           => n529, outb => n747);
   U939 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_1_0_port, b
                           => n530, c => 
                           load_n_store_RGB_Array_2_block_ram_r_0_0_port, d => 
                           n531, outb => n746);
   U940 : aoi22 port map( a => n532, b => n686, c => n534, d => n704, outb => 
                           n744);
   U941 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_2_0_port, 
                           outb => n704);
   U942 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_4_0_port, 
                           outb => n686);
   U943 : nand2 port map( a => n536, b => n668, outb => n743);
   U944 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_6_0_port, 
                           outb => n668);
   U945 : nand4 port map( a => n538, b => n749, c => n750, d => n751, outb => 
                           n740);
   U946 : nor3 port map( a => n752, b => n753, c => n754, outb => n751);
   U947 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_13_0_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_2_block_ram_r_11_0_port, d =>
                           n528, outb => n754);
   U948 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_15_0_port, b
                           => n529, outb => n753);
   U949 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_9_0_port, b
                           => n530, c => 
                           load_n_store_RGB_Array_2_block_ram_r_8_0_port, d => 
                           n531, outb => n752);
   U950 : aoi22 port map( a => n532, b => n612, c => n534, d => n630, outb => 
                           n750);
   U951 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_10_0_port, 
                           outb => n630);
   U952 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_12_0_port, 
                           outb => n612);
   U953 : nand2 port map( a => n536, b => n594, outb => n749);
   U954 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_14_0_port, 
                           outb => n594);
   U955 : nand3 port map( a => n755, b => n756, c => n757, outb => n2308);
   U956 : nand2 port map( a => load_n_store_lazy_in_2_7_port, b => 
                           load_n_store_we_i, outb => n757);
   U957 : nand4 port map( a => n520, b => n758, c => n759, d => n760, outb => 
                           n756);
   U958 : nor3 port map( a => n761, b => n762, c => n763, outb => n760);
   U959 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_5_7_port, b
                           => n527, c => 
                           load_n_store_RGB_Array_2_block_ram_r_3_7_port, d => 
                           n528, outb => n763);
   U960 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_7_7_port, b 
                           => n529, outb => n762);
   U961 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_1_7_port, b
                           => n530, c => 
                           load_n_store_RGB_Array_2_block_ram_r_0_7_port, d => 
                           n531, outb => n761);
   U962 : aoi22 port map( a => n532, b => n681, c => n534, d => n699, outb => 
                           n759);
   U963 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_2_7_port, 
                           outb => n699);
   U964 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_4_7_port, 
                           outb => n681);
   U965 : nand2 port map( a => n536, b => n663, outb => n758);
   U966 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_6_7_port, 
                           outb => n663);
   U967 : nand4 port map( a => n538, b => n764, c => n765, d => n766, outb => 
                           n755);
   U968 : nor3 port map( a => n767, b => n768, c => n769, outb => n766);
   U969 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_13_7_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_2_block_ram_r_11_7_port, d =>
                           n528, outb => n769);
   U970 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_15_7_port, b
                           => n529, outb => n768);
   U971 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_9_7_port, b
                           => n530, c => 
                           load_n_store_RGB_Array_2_block_ram_r_8_7_port, d => 
                           n531, outb => n767);
   U972 : aoi22 port map( a => n532, b => n607, c => n534, d => n625, outb => 
                           n765);
   U973 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_10_7_port, 
                           outb => n625);
   U974 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_12_7_port, 
                           outb => n607);
   U975 : nand2 port map( a => n536, b => n561, outb => n764);
   U976 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_14_7_port, 
                           outb => n561);
   U977 : nand3 port map( a => n770, b => n771, c => n772, outb => n2307);
   U978 : nand2 port map( a => load_n_store_lazy_in_2_6_port, b => 
                           load_n_store_we_i, outb => n772);
   U979 : nand4 port map( a => n520, b => n773, c => n774, d => n775, outb => 
                           n771);
   U980 : nor3 port map( a => n776, b => n777, c => n778, outb => n775);
   U981 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_5_6_port, b
                           => n527, c => 
                           load_n_store_RGB_Array_2_block_ram_r_3_6_port, d => 
                           n528, outb => n778);
   U982 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_7_6_port, b 
                           => n529, outb => n777);
   U983 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_1_6_port, b
                           => n530, c => 
                           load_n_store_RGB_Array_2_block_ram_r_0_6_port, d => 
                           n531, outb => n776);
   U984 : aoi22 port map( a => n532, b => n682, c => n534, d => n700, outb => 
                           n774);
   U985 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_2_6_port, 
                           outb => n700);
   U986 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_4_6_port, 
                           outb => n682);
   U987 : nand2 port map( a => n536, b => n664, outb => n773);
   U988 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_6_6_port, 
                           outb => n664);
   U989 : nand4 port map( a => n538, b => n779, c => n780, d => n781, outb => 
                           n770);
   U990 : nor3 port map( a => n782, b => n783, c => n784, outb => n781);
   U991 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_13_6_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_2_block_ram_r_11_6_port, d =>
                           n528, outb => n784);
   U992 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_15_6_port, b
                           => n529, outb => n783);
   U993 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_9_6_port, b
                           => n530, c => 
                           load_n_store_RGB_Array_2_block_ram_r_8_6_port, d => 
                           n531, outb => n782);
   U994 : aoi22 port map( a => n532, b => n608, c => n534, d => n626, outb => 
                           n780);
   U995 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_10_6_port, 
                           outb => n626);
   U996 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_12_6_port, 
                           outb => n608);
   U997 : nand2 port map( a => n536, b => n563, outb => n779);
   U998 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_14_6_port, 
                           outb => n563);
   U999 : nand3 port map( a => n785, b => n786, c => n787, outb => n2306);
   U1000 : nand2 port map( a => load_n_store_lazy_in_2_5_port, b => 
                           load_n_store_we_i, outb => n787);
   U1001 : nand4 port map( a => n520, b => n788, c => n789, d => n790, outb => 
                           n786);
   U1002 : nor3 port map( a => n791, b => n792, c => n793, outb => n790);
   U1003 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_5_5_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_2_block_ram_r_3_5_port, d => 
                           n528, outb => n793);
   U1004 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_7_5_port, b
                           => n529, outb => n792);
   U1005 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_1_5_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_2_block_ram_r_0_5_port, d => 
                           n531, outb => n791);
   U1006 : aoi22 port map( a => n532, b => n683, c => n534, d => n701, outb => 
                           n789);
   U1007 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_2_5_port, 
                           outb => n701);
   U1008 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_4_5_port, 
                           outb => n683);
   U1009 : nand2 port map( a => n536, b => n665, outb => n788);
   U1010 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_6_5_port, 
                           outb => n665);
   U1011 : nand4 port map( a => n538, b => n794, c => n795, d => n796, outb => 
                           n785);
   U1012 : nor3 port map( a => n797, b => n798, c => n799, outb => n796);
   U1013 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_13_5_port,
                           b => n527, c => 
                           load_n_store_RGB_Array_2_block_ram_r_11_5_port, d =>
                           n528, outb => n799);
   U1014 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_15_5_port, 
                           b => n529, outb => n798);
   U1015 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_9_5_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_2_block_ram_r_8_5_port, d => 
                           n531, outb => n797);
   U1016 : aoi22 port map( a => n532, b => n609, c => n534, d => n627, outb => 
                           n795);
   U1017 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_10_5_port,
                           outb => n627);
   U1018 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_12_5_port,
                           outb => n609);
   U1019 : nand2 port map( a => n536, b => n565, outb => n794);
   U1020 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_14_5_port,
                           outb => n565);
   U1021 : nand3 port map( a => n800, b => n801, c => n802, outb => n2305);
   U1022 : nand2 port map( a => load_n_store_lazy_in_2_4_port, b => 
                           load_n_store_we_i, outb => n802);
   U1023 : nand4 port map( a => n520, b => n803, c => n804, d => n805, outb => 
                           n801);
   U1024 : nor3 port map( a => n806, b => n807, c => n808, outb => n805);
   U1025 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_5_4_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_2_block_ram_r_3_4_port, d => 
                           n528, outb => n808);
   U1026 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_7_4_port, b
                           => n529, outb => n807);
   U1027 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_1_4_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_2_block_ram_r_0_4_port, d => 
                           n531, outb => n806);
   U1028 : aoi22 port map( a => n532, b => n684, c => n534, d => n702, outb => 
                           n804);
   U1029 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_2_4_port, 
                           outb => n702);
   U1030 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_4_4_port, 
                           outb => n684);
   U1031 : nand2 port map( a => n536, b => n666, outb => n803);
   U1032 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_6_4_port, 
                           outb => n666);
   U1033 : nand4 port map( a => n538, b => n809, c => n810, d => n811, outb => 
                           n800);
   U1034 : nor3 port map( a => n812, b => n813, c => n814, outb => n811);
   U1035 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_13_4_port,
                           b => n527, c => 
                           load_n_store_RGB_Array_2_block_ram_r_11_4_port, d =>
                           n528, outb => n814);
   U1036 : nor2 port map( a => load_n_store_RGB_Array_2_block_ram_r_15_4_port, 
                           b => n529, outb => n813);
   U1037 : oai22 port map( a => load_n_store_RGB_Array_2_block_ram_r_9_4_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_2_block_ram_r_8_4_port, d => 
                           n531, outb => n812);
   U1038 : aoi22 port map( a => n532, b => n610, c => n534, d => n628, outb => 
                           n810);
   U1039 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_10_4_port,
                           outb => n628);
   U1040 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_12_4_port,
                           outb => n610);
   U1041 : nand2 port map( a => n536, b => n588, outb => n809);
   U1042 : inv port map( inb => load_n_store_RGB_Array_2_block_ram_r_14_4_port,
                           outb => n588);
   U1043 : nand3 port map( a => n815, b => n816, c => n817, outb => n2032);
   U1044 : nand2 port map( a => load_n_store_lazy_in_1_3_port, b => 
                           load_n_store_we_i, outb => n817);
   U1045 : nand4 port map( a => n520, b => n818, c => n819, d => n820, outb => 
                           n816);
   U1046 : nor3 port map( a => n821, b => n822, c => n823, outb => n820);
   U1047 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_5_3_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_1_block_ram_r_3_3_port, d => 
                           n528, outb => n823);
   U1048 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_7_3_port, b
                           => n529, outb => n822);
   U1049 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_1_3_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_1_block_ram_r_0_3_port, d => 
                           n531, outb => n821);
   U1050 : aoi22 port map( a => n532, b => n824, c => n534, d => n825, outb => 
                           n819);
   U1051 : nand2 port map( a => n536, b => n826, outb => n818);
   U1052 : nand4 port map( a => n538, b => n827, c => n828, d => n829, outb => 
                           n815);
   U1053 : nor3 port map( a => n830, b => n831, c => n832, outb => n829);
   U1054 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_13_3_port,
                           b => n527, c => 
                           load_n_store_RGB_Array_1_block_ram_r_11_3_port, d =>
                           n528, outb => n832);
   U1055 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_15_3_port, 
                           b => n529, outb => n831);
   U1056 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_9_3_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_1_block_ram_r_8_3_port, d => 
                           n531, outb => n830);
   U1057 : aoi22 port map( a => n532, b => n833, c => n534, d => n834, outb => 
                           n828);
   U1058 : nand2 port map( a => n536, b => n835, outb => n827);
   U1059 : inv port map( inb => n836, outb => n2300);
   U1060 : aoi22 port map( a => load_n_store_lazy_in_1_7_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_1_block_ram_r_15_7_port, outb
                           => n836);
   U1061 : inv port map( inb => n837, outb => n2299);
   U1062 : aoi22 port map( a => load_n_store_lazy_in_1_6_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_1_block_ram_r_15_6_port, outb
                           => n837);
   U1063 : inv port map( inb => n838, outb => n2298);
   U1064 : aoi22 port map( a => load_n_store_lazy_in_1_5_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_1_block_ram_r_15_5_port, outb
                           => n838);
   U1065 : inv port map( inb => n839, outb => n2297);
   U1066 : aoi22 port map( a => load_n_store_lazy_in_1_4_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_1_block_ram_r_15_4_port, outb
                           => n839);
   U1067 : inv port map( inb => n840, outb => n2296);
   U1068 : aoi22 port map( a => load_n_store_lazy_in_1_3_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_1_block_ram_r_15_3_port, outb
                           => n840);
   U1069 : inv port map( inb => n841, outb => n2295);
   U1070 : aoi22 port map( a => load_n_store_lazy_in_1_2_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_1_block_ram_r_15_2_port, outb
                           => n841);
   U1071 : inv port map( inb => n842, outb => n2294);
   U1072 : aoi22 port map( a => load_n_store_lazy_in_1_1_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_1_block_ram_r_15_1_port, outb
                           => n842);
   U1073 : inv port map( inb => n843, outb => n2293);
   U1074 : aoi22 port map( a => load_n_store_lazy_in_1_0_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_1_block_ram_r_15_0_port, outb
                           => n843);
   U1075 : oai22 port map( a => n844, b => n559, c => n560, d => n845, outb => 
                           n2292);
   U1076 : oai22 port map( a => n846, b => n559, c => n560, d => n847, outb => 
                           n2291);
   U1077 : oai22 port map( a => n848, b => n559, c => n560, d => n849, outb => 
                           n2290);
   U1078 : nand3 port map( a => n850, b => n851, c => n852, outb => n2031);
   U1079 : nand2 port map( a => load_n_store_lazy_in_1_2_port, b => 
                           load_n_store_we_i, outb => n852);
   U1080 : nand4 port map( a => n520, b => n853, c => n854, d => n855, outb => 
                           n851);
   U1081 : nor3 port map( a => n856, b => n857, c => n858, outb => n855);
   U1082 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_5_2_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_1_block_ram_r_3_2_port, d => 
                           n528, outb => n858);
   U1083 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_7_2_port, b
                           => n529, outb => n857);
   U1084 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_1_2_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_1_block_ram_r_0_2_port, d => 
                           n531, outb => n856);
   U1085 : aoi22 port map( a => n532, b => n859, c => n534, d => n860, outb => 
                           n854);
   U1086 : nand2 port map( a => n536, b => n861, outb => n853);
   U1087 : nand4 port map( a => n538, b => n862, c => n863, d => n864, outb => 
                           n850);
   U1088 : nor3 port map( a => n865, b => n866, c => n867, outb => n864);
   U1089 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_13_2_port,
                           b => n527, c => 
                           load_n_store_RGB_Array_1_block_ram_r_11_2_port, d =>
                           n528, outb => n867);
   U1090 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_15_2_port, 
                           b => n529, outb => n866);
   U1091 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_9_2_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_1_block_ram_r_8_2_port, d => 
                           n531, outb => n865);
   U1092 : aoi22 port map( a => n532, b => n868, c => n534, d => n869, outb => 
                           n863);
   U1093 : nand2 port map( a => n536, b => n870, outb => n862);
   U1094 : oai22 port map( a => n871, b => n559, c => n560, d => n872, outb => 
                           n2289);
   U1095 : oai22 port map( a => n873, b => n559, c => n560, d => n835, outb => 
                           n2288);
   U1096 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_14_3_port,
                           outb => n835);
   U1097 : oai22 port map( a => n874, b => n559, c => n560, d => n870, outb => 
                           n2287);
   U1098 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_14_2_port,
                           outb => n870);
   U1099 : oai22 port map( a => n875, b => n559, c => n560, d => n876, outb => 
                           n2286);
   U1100 : oai22 port map( a => n877, b => n559, c => n560, d => n878, outb => 
                           n2285);
   U1101 : inv port map( inb => n879, outb => n2284);
   U1102 : aoi22 port map( a => load_n_store_lazy_in_1_7_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_1_block_ram_r_13_7_port, outb
                           => n879);
   U1103 : inv port map( inb => n880, outb => n2283);
   U1104 : aoi22 port map( a => load_n_store_lazy_in_1_6_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_1_block_ram_r_13_6_port, outb
                           => n880);
   U1105 : inv port map( inb => n881, outb => n2282);
   U1106 : aoi22 port map( a => load_n_store_lazy_in_1_5_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_1_block_ram_r_13_5_port, outb
                           => n881);
   U1107 : inv port map( inb => n882, outb => n2281);
   U1108 : aoi22 port map( a => load_n_store_lazy_in_1_4_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_1_block_ram_r_13_4_port, outb
                           => n882);
   U1109 : inv port map( inb => n883, outb => n2280);
   U1110 : aoi22 port map( a => load_n_store_lazy_in_1_3_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_1_block_ram_r_13_3_port, outb
                           => n883);
   U1111 : inv port map( inb => n884, outb => n2279);
   U1112 : aoi22 port map( a => load_n_store_lazy_in_1_2_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_1_block_ram_r_13_2_port, outb
                           => n884);
   U1113 : inv port map( inb => n885, outb => n2278);
   U1114 : aoi22 port map( a => load_n_store_lazy_in_1_1_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_1_block_ram_r_13_1_port, outb
                           => n885);
   U1115 : inv port map( inb => n886, outb => n2277);
   U1116 : aoi22 port map( a => load_n_store_lazy_in_1_0_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_1_block_ram_r_13_0_port, outb
                           => n886);
   U1117 : oai22 port map( a => n844, b => n605, c => n606, d => n887, outb => 
                           n2276);
   U1118 : oai22 port map( a => n846, b => n605, c => n606, d => n888, outb => 
                           n2275);
   U1119 : oai22 port map( a => n848, b => n605, c => n606, d => n889, outb => 
                           n2274);
   U1120 : oai22 port map( a => n871, b => n605, c => n606, d => n890, outb => 
                           n2273);
   U1121 : oai22 port map( a => n873, b => n605, c => n606, d => n833, outb => 
                           n2272);
   U1122 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_12_3_port,
                           outb => n833);
   U1123 : oai22 port map( a => n874, b => n605, c => n606, d => n868, outb => 
                           n2271);
   U1124 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_12_2_port,
                           outb => n868);
   U1125 : oai22 port map( a => n875, b => n605, c => n606, d => n891, outb => 
                           n2270);
   U1126 : oai22 port map( a => n877, b => n605, c => n606, d => n892, outb => 
                           n2269);
   U1127 : inv port map( inb => n893, outb => n2268);
   U1128 : aoi22 port map( a => load_n_store_lazy_in_1_7_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_1_block_ram_r_11_7_port, outb
                           => n893);
   U1129 : inv port map( inb => n894, outb => n2267);
   U1130 : aoi22 port map( a => load_n_store_lazy_in_1_6_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_1_block_ram_r_11_6_port, outb
                           => n894);
   U1131 : inv port map( inb => n895, outb => n2266);
   U1132 : aoi22 port map( a => load_n_store_lazy_in_1_5_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_1_block_ram_r_11_5_port, outb
                           => n895);
   U1133 : inv port map( inb => n896, outb => n2265);
   U1134 : aoi22 port map( a => load_n_store_lazy_in_1_4_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_1_block_ram_r_11_4_port, outb
                           => n896);
   U1135 : inv port map( inb => n897, outb => n2264);
   U1136 : aoi22 port map( a => load_n_store_lazy_in_1_3_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_1_block_ram_r_11_3_port, outb
                           => n897);
   U1137 : inv port map( inb => n898, outb => n2263);
   U1138 : aoi22 port map( a => load_n_store_lazy_in_1_2_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_1_block_ram_r_11_2_port, outb
                           => n898);
   U1139 : inv port map( inb => n899, outb => n2262);
   U1140 : aoi22 port map( a => load_n_store_lazy_in_1_1_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_1_block_ram_r_11_1_port, outb
                           => n899);
   U1141 : inv port map( inb => n900, outb => n2261);
   U1142 : aoi22 port map( a => load_n_store_lazy_in_1_0_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_1_block_ram_r_11_0_port, outb
                           => n900);
   U1143 : oai22 port map( a => n844, b => n623, c => n624, d => n901, outb => 
                           n2260);
   U1144 : oai22 port map( a => n846, b => n623, c => n624, d => n902, outb => 
                           n2259);
   U1145 : oai22 port map( a => n848, b => n623, c => n624, d => n903, outb => 
                           n2258);
   U1146 : oai22 port map( a => n871, b => n623, c => n624, d => n904, outb => 
                           n2257);
   U1147 : oai22 port map( a => n873, b => n623, c => n624, d => n834, outb => 
                           n2256);
   U1148 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_10_3_port,
                           outb => n834);
   U1149 : oai22 port map( a => n874, b => n623, c => n624, d => n869, outb => 
                           n2255);
   U1150 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_10_2_port,
                           outb => n869);
   U1151 : oai22 port map( a => n875, b => n623, c => n624, d => n905, outb => 
                           n2254);
   U1152 : oai22 port map( a => n877, b => n623, c => n624, d => n906, outb => 
                           n2253);
   U1153 : inv port map( inb => n907, outb => n2252);
   U1154 : aoi22 port map( a => load_n_store_lazy_in_1_7_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_1_block_ram_r_9_7_port, outb 
                           => n907);
   U1155 : inv port map( inb => n908, outb => n2251);
   U1156 : aoi22 port map( a => load_n_store_lazy_in_1_6_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_1_block_ram_r_9_6_port, outb 
                           => n908);
   U1157 : inv port map( inb => n909, outb => n2250);
   U1158 : aoi22 port map( a => load_n_store_lazy_in_1_5_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_1_block_ram_r_9_5_port, outb 
                           => n909);
   U1159 : inv port map( inb => n910, outb => n2249);
   U1160 : aoi22 port map( a => load_n_store_lazy_in_1_4_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_1_block_ram_r_9_4_port, outb 
                           => n910);
   U1161 : inv port map( inb => n911, outb => n2248);
   U1162 : aoi22 port map( a => load_n_store_lazy_in_1_3_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_1_block_ram_r_9_3_port, outb 
                           => n911);
   U1163 : inv port map( inb => n912, outb => n2247);
   U1164 : aoi22 port map( a => load_n_store_lazy_in_1_2_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_1_block_ram_r_9_2_port, outb 
                           => n912);
   U1165 : inv port map( inb => n913, outb => n2246);
   U1166 : aoi22 port map( a => load_n_store_lazy_in_1_1_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_1_block_ram_r_9_1_port, outb 
                           => n913);
   U1167 : inv port map( inb => n914, outb => n2245);
   U1168 : aoi22 port map( a => load_n_store_lazy_in_1_0_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_1_block_ram_r_9_0_port, outb 
                           => n914);
   U1169 : inv port map( inb => n915, outb => n2244);
   U1170 : aoi22 port map( a => load_n_store_lazy_in_1_7_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_1_block_ram_r_8_7_port, outb 
                           => n915);
   U1171 : inv port map( inb => n916, outb => n2243);
   U1172 : aoi22 port map( a => load_n_store_lazy_in_1_6_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_1_block_ram_r_8_6_port, outb 
                           => n916);
   U1173 : inv port map( inb => n917, outb => n2242);
   U1174 : aoi22 port map( a => load_n_store_lazy_in_1_5_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_1_block_ram_r_8_5_port, outb 
                           => n917);
   U1175 : inv port map( inb => n918, outb => n2241);
   U1176 : aoi22 port map( a => load_n_store_lazy_in_1_4_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_1_block_ram_r_8_4_port, outb 
                           => n918);
   U1177 : inv port map( inb => n919, outb => n2240);
   U1178 : aoi22 port map( a => load_n_store_lazy_in_1_3_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_1_block_ram_r_8_3_port, outb 
                           => n919);
   U1179 : inv port map( inb => n920, outb => n2239);
   U1180 : aoi22 port map( a => load_n_store_lazy_in_1_2_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_1_block_ram_r_8_2_port, outb 
                           => n920);
   U1181 : inv port map( inb => n921, outb => n2238);
   U1182 : aoi22 port map( a => load_n_store_lazy_in_1_1_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_1_block_ram_r_8_1_port, outb 
                           => n921);
   U1183 : inv port map( inb => n922, outb => n2237);
   U1184 : aoi22 port map( a => load_n_store_lazy_in_1_0_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_1_block_ram_r_8_0_port, outb 
                           => n922);
   U1185 : inv port map( inb => n923, outb => n2236);
   U1186 : aoi22 port map( a => load_n_store_lazy_in_1_7_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_1_block_ram_r_7_7_port, outb 
                           => n923);
   U1187 : inv port map( inb => n924, outb => n2235);
   U1188 : aoi22 port map( a => load_n_store_lazy_in_1_6_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_1_block_ram_r_7_6_port, outb 
                           => n924);
   U1189 : inv port map( inb => n925, outb => n2234);
   U1190 : aoi22 port map( a => load_n_store_lazy_in_1_5_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_1_block_ram_r_7_5_port, outb 
                           => n925);
   U1191 : inv port map( inb => n926, outb => n2233);
   U1192 : aoi22 port map( a => load_n_store_lazy_in_1_4_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_1_block_ram_r_7_4_port, outb 
                           => n926);
   U1193 : inv port map( inb => n927, outb => n2232);
   U1194 : aoi22 port map( a => load_n_store_lazy_in_1_3_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_1_block_ram_r_7_3_port, outb 
                           => n927);
   U1195 : inv port map( inb => n928, outb => n2231);
   U1196 : aoi22 port map( a => load_n_store_lazy_in_1_2_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_1_block_ram_r_7_2_port, outb 
                           => n928);
   U1197 : inv port map( inb => n929, outb => n2230);
   U1198 : aoi22 port map( a => load_n_store_lazy_in_1_1_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_1_block_ram_r_7_1_port, outb 
                           => n929);
   U1199 : inv port map( inb => n930, outb => n2229);
   U1200 : aoi22 port map( a => load_n_store_lazy_in_1_0_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_1_block_ram_r_7_0_port, outb 
                           => n930);
   U1201 : oai22 port map( a => n844, b => n661, c => n662, d => n931, outb => 
                           n2228);
   U1202 : oai22 port map( a => n846, b => n661, c => n662, d => n932, outb => 
                           n2227);
   U1203 : oai22 port map( a => n848, b => n661, c => n662, d => n933, outb => 
                           n2226);
   U1204 : oai22 port map( a => n871, b => n661, c => n662, d => n934, outb => 
                           n2225);
   U1205 : oai22 port map( a => n873, b => n661, c => n662, d => n826, outb => 
                           n2224);
   U1206 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_6_3_port, 
                           outb => n826);
   U1207 : oai22 port map( a => n874, b => n661, c => n662, d => n861, outb => 
                           n2223);
   U1208 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_6_2_port, 
                           outb => n861);
   U1209 : oai22 port map( a => n875, b => n661, c => n662, d => n935, outb => 
                           n2222);
   U1210 : oai22 port map( a => n877, b => n661, c => n662, d => n936, outb => 
                           n2221);
   U1211 : inv port map( inb => n937, outb => n2220);
   U1212 : aoi22 port map( a => load_n_store_lazy_in_1_7_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_1_block_ram_r_5_7_port, outb 
                           => n937);
   U1213 : inv port map( inb => n938, outb => n2219);
   U1214 : aoi22 port map( a => load_n_store_lazy_in_1_6_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_1_block_ram_r_5_6_port, outb 
                           => n938);
   U1215 : inv port map( inb => n939, outb => n2218);
   U1216 : aoi22 port map( a => load_n_store_lazy_in_1_5_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_1_block_ram_r_5_5_port, outb 
                           => n939);
   U1217 : inv port map( inb => n940, outb => n2217);
   U1218 : aoi22 port map( a => load_n_store_lazy_in_1_4_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_1_block_ram_r_5_4_port, outb 
                           => n940);
   U1219 : inv port map( inb => n941, outb => n2216);
   U1220 : aoi22 port map( a => load_n_store_lazy_in_1_3_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_1_block_ram_r_5_3_port, outb 
                           => n941);
   U1221 : inv port map( inb => n942, outb => n2215);
   U1222 : aoi22 port map( a => load_n_store_lazy_in_1_2_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_1_block_ram_r_5_2_port, outb 
                           => n942);
   U1223 : inv port map( inb => n943, outb => n2214);
   U1224 : aoi22 port map( a => load_n_store_lazy_in_1_1_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_1_block_ram_r_5_1_port, outb 
                           => n943);
   U1225 : inv port map( inb => n944, outb => n2213);
   U1226 : aoi22 port map( a => load_n_store_lazy_in_1_0_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_1_block_ram_r_5_0_port, outb 
                           => n944);
   U1227 : oai22 port map( a => n844, b => n679, c => n680, d => n945, outb => 
                           n2212);
   U1228 : oai22 port map( a => n846, b => n679, c => n680, d => n946, outb => 
                           n2211);
   U1229 : oai22 port map( a => n848, b => n679, c => n680, d => n947, outb => 
                           n2210);
   U1230 : oai22 port map( a => n871, b => n679, c => n680, d => n948, outb => 
                           n2209);
   U1231 : oai22 port map( a => n873, b => n679, c => n680, d => n824, outb => 
                           n2208);
   U1232 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_4_3_port, 
                           outb => n824);
   U1233 : oai22 port map( a => n874, b => n679, c => n680, d => n859, outb => 
                           n2207);
   U1234 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_4_2_port, 
                           outb => n859);
   U1235 : oai22 port map( a => n875, b => n679, c => n680, d => n949, outb => 
                           n2206);
   U1236 : oai22 port map( a => n877, b => n679, c => n680, d => n950, outb => 
                           n2205);
   U1237 : inv port map( inb => n951, outb => n2204);
   U1238 : aoi22 port map( a => load_n_store_lazy_in_1_7_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_1_block_ram_r_3_7_port, outb 
                           => n951);
   U1239 : inv port map( inb => n952, outb => n2203);
   U1240 : aoi22 port map( a => load_n_store_lazy_in_1_6_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_1_block_ram_r_3_6_port, outb 
                           => n952);
   U1241 : inv port map( inb => n953, outb => n2202);
   U1242 : aoi22 port map( a => load_n_store_lazy_in_1_5_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_1_block_ram_r_3_5_port, outb 
                           => n953);
   U1243 : inv port map( inb => n954, outb => n2201);
   U1244 : aoi22 port map( a => load_n_store_lazy_in_1_4_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_1_block_ram_r_3_4_port, outb 
                           => n954);
   U1245 : inv port map( inb => n955, outb => n2200);
   U1246 : aoi22 port map( a => load_n_store_lazy_in_1_3_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_1_block_ram_r_3_3_port, outb 
                           => n955);
   U1247 : inv port map( inb => n956, outb => n2199);
   U1248 : aoi22 port map( a => load_n_store_lazy_in_1_2_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_1_block_ram_r_3_2_port, outb 
                           => n956);
   U1249 : inv port map( inb => n957, outb => n2198);
   U1250 : aoi22 port map( a => load_n_store_lazy_in_1_1_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_1_block_ram_r_3_1_port, outb 
                           => n957);
   U1251 : inv port map( inb => n958, outb => n2197);
   U1252 : aoi22 port map( a => load_n_store_lazy_in_1_0_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_1_block_ram_r_3_0_port, outb 
                           => n958);
   U1253 : oai22 port map( a => n844, b => n697, c => n698, d => n959, outb => 
                           n2196);
   U1254 : inv port map( inb => load_n_store_lazy_in_1_7_port, outb => n844);
   U1255 : oai22 port map( a => n846, b => n697, c => n698, d => n960, outb => 
                           n2195);
   U1256 : inv port map( inb => load_n_store_lazy_in_1_6_port, outb => n846);
   U1257 : oai22 port map( a => n848, b => n697, c => n698, d => n961, outb => 
                           n2194);
   U1258 : inv port map( inb => load_n_store_lazy_in_1_5_port, outb => n848);
   U1259 : oai22 port map( a => n871, b => n697, c => n698, d => n962, outb => 
                           n2193);
   U1260 : inv port map( inb => load_n_store_lazy_in_1_4_port, outb => n871);
   U1261 : oai22 port map( a => n873, b => n697, c => n698, d => n825, outb => 
                           n2192);
   U1262 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_2_3_port, 
                           outb => n825);
   U1263 : inv port map( inb => load_n_store_lazy_in_1_3_port, outb => n873);
   U1264 : oai22 port map( a => n874, b => n697, c => n698, d => n860, outb => 
                           n2191);
   U1265 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_2_2_port, 
                           outb => n860);
   U1266 : inv port map( inb => load_n_store_lazy_in_1_2_port, outb => n874);
   U1267 : oai22 port map( a => n875, b => n697, c => n698, d => n963, outb => 
                           n2190);
   U1268 : inv port map( inb => load_n_store_lazy_in_1_1_port, outb => n875);
   U1269 : oai22 port map( a => n877, b => n697, c => n698, d => n964, outb => 
                           n2189);
   U1270 : inv port map( inb => load_n_store_lazy_in_1_0_port, outb => n877);
   U1271 : inv port map( inb => n965, outb => n2188);
   U1272 : aoi22 port map( a => load_n_store_lazy_in_1_7_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_1_block_ram_r_1_7_port, outb 
                           => n965);
   U1273 : inv port map( inb => n966, outb => n2187);
   U1274 : aoi22 port map( a => load_n_store_lazy_in_1_6_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_1_block_ram_r_1_6_port, outb 
                           => n966);
   U1275 : inv port map( inb => n967, outb => n2186);
   U1276 : aoi22 port map( a => load_n_store_lazy_in_1_5_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_1_block_ram_r_1_5_port, outb 
                           => n967);
   U1277 : inv port map( inb => n968, outb => n2185);
   U1278 : aoi22 port map( a => load_n_store_lazy_in_1_4_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_1_block_ram_r_1_4_port, outb 
                           => n968);
   U1279 : inv port map( inb => n969, outb => n2184);
   U1280 : aoi22 port map( a => load_n_store_lazy_in_1_3_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_1_block_ram_r_1_3_port, outb 
                           => n969);
   U1281 : inv port map( inb => n970, outb => n2183);
   U1282 : aoi22 port map( a => load_n_store_lazy_in_1_2_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_1_block_ram_r_1_2_port, outb 
                           => n970);
   U1283 : inv port map( inb => n971, outb => n2182);
   U1284 : aoi22 port map( a => load_n_store_lazy_in_1_1_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_1_block_ram_r_1_1_port, outb 
                           => n971);
   U1285 : inv port map( inb => n972, outb => n2181);
   U1286 : aoi22 port map( a => load_n_store_lazy_in_1_0_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_1_block_ram_r_1_0_port, outb 
                           => n972);
   U1287 : inv port map( inb => n973, outb => n2180);
   U1288 : aoi22 port map( a => load_n_store_lazy_in_1_7_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_1_block_ram_r_0_7_port, outb 
                           => n973);
   U1289 : inv port map( inb => n974, outb => n2179);
   U1290 : aoi22 port map( a => load_n_store_lazy_in_1_6_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_1_block_ram_r_0_6_port, outb 
                           => n974);
   U1291 : inv port map( inb => n975, outb => n2178);
   U1292 : aoi22 port map( a => load_n_store_lazy_in_1_5_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_1_block_ram_r_0_5_port, outb 
                           => n975);
   U1293 : inv port map( inb => n976, outb => n2177);
   U1294 : aoi22 port map( a => load_n_store_lazy_in_1_4_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_1_block_ram_r_0_4_port, outb 
                           => n976);
   U1295 : inv port map( inb => n977, outb => n2176);
   U1296 : aoi22 port map( a => load_n_store_lazy_in_1_3_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_1_block_ram_r_0_3_port, outb 
                           => n977);
   U1297 : inv port map( inb => n978, outb => n2175);
   U1298 : aoi22 port map( a => load_n_store_lazy_in_1_2_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_1_block_ram_r_0_2_port, outb 
                           => n978);
   U1299 : inv port map( inb => n979, outb => n2174);
   U1300 : aoi22 port map( a => load_n_store_lazy_in_1_1_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_1_block_ram_r_0_1_port, outb 
                           => n979);
   U1301 : inv port map( inb => n980, outb => n2173);
   U1302 : aoi22 port map( a => load_n_store_lazy_in_1_0_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_1_block_ram_r_0_0_port, outb 
                           => n980);
   U1303 : nand3 port map( a => n981, b => n982, c => n983, outb => n2030);
   U1304 : nand2 port map( a => load_n_store_lazy_in_1_1_port, b => 
                           load_n_store_we_i, outb => n983);
   U1305 : nand4 port map( a => n520, b => n984, c => n985, d => n986, outb => 
                           n982);
   U1306 : nor3 port map( a => n987, b => n988, c => n989, outb => n986);
   U1307 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_5_1_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_1_block_ram_r_3_1_port, d => 
                           n528, outb => n989);
   U1308 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_7_1_port, b
                           => n529, outb => n988);
   U1309 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_1_1_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_1_block_ram_r_0_1_port, d => 
                           n531, outb => n987);
   U1310 : aoi22 port map( a => n532, b => n949, c => n534, d => n963, outb => 
                           n985);
   U1311 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_2_1_port, 
                           outb => n963);
   U1312 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_4_1_port, 
                           outb => n949);
   U1313 : nand2 port map( a => n536, b => n935, outb => n984);
   U1314 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_6_1_port, 
                           outb => n935);
   U1315 : nand4 port map( a => n538, b => n990, c => n991, d => n992, outb => 
                           n981);
   U1316 : nor3 port map( a => n993, b => n994, c => n995, outb => n992);
   U1317 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_13_1_port,
                           b => n527, c => 
                           load_n_store_RGB_Array_1_block_ram_r_11_1_port, d =>
                           n528, outb => n995);
   U1318 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_15_1_port, 
                           b => n529, outb => n994);
   U1319 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_9_1_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_1_block_ram_r_8_1_port, d => 
                           n531, outb => n993);
   U1320 : aoi22 port map( a => n532, b => n891, c => n534, d => n905, outb => 
                           n991);
   U1321 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_10_1_port,
                           outb => n905);
   U1322 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_12_1_port,
                           outb => n891);
   U1323 : nand2 port map( a => n536, b => n876, outb => n990);
   U1324 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_14_1_port,
                           outb => n876);
   U1325 : nand3 port map( a => n996, b => n997, c => n998, outb => n2029);
   U1326 : nand2 port map( a => load_n_store_lazy_in_1_0_port, b => 
                           load_n_store_we_i, outb => n998);
   U1327 : nand4 port map( a => n520, b => n999, c => n1000, d => n1001, outb 
                           => n997);
   U1328 : nor3 port map( a => n1002, b => n1003, c => n1004, outb => n1001);
   U1329 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_5_0_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_1_block_ram_r_3_0_port, d => 
                           n528, outb => n1004);
   U1330 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_7_0_port, b
                           => n529, outb => n1003);
   U1331 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_1_0_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_1_block_ram_r_0_0_port, d => 
                           n531, outb => n1002);
   U1332 : aoi22 port map( a => n532, b => n950, c => n534, d => n964, outb => 
                           n1000);
   U1333 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_2_0_port, 
                           outb => n964);
   U1334 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_4_0_port, 
                           outb => n950);
   U1335 : nand2 port map( a => n536, b => n936, outb => n999);
   U1336 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_6_0_port, 
                           outb => n936);
   U1337 : nand4 port map( a => n538, b => n1005, c => n1006, d => n1007, outb 
                           => n996);
   U1338 : nor3 port map( a => n1008, b => n1009, c => n1010, outb => n1007);
   U1339 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_13_0_port,
                           b => n527, c => 
                           load_n_store_RGB_Array_1_block_ram_r_11_0_port, d =>
                           n528, outb => n1010);
   U1340 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_15_0_port, 
                           b => n529, outb => n1009);
   U1341 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_9_0_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_1_block_ram_r_8_0_port, d => 
                           n531, outb => n1008);
   U1342 : aoi22 port map( a => n532, b => n892, c => n534, d => n906, outb => 
                           n1006);
   U1343 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_10_0_port,
                           outb => n906);
   U1344 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_12_0_port,
                           outb => n892);
   U1345 : nand2 port map( a => n536, b => n878, outb => n1005);
   U1346 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_14_0_port,
                           outb => n878);
   U1347 : nand3 port map( a => n1011, b => n1012, c => n1013, outb => n2036);
   U1348 : nand2 port map( a => load_n_store_lazy_in_1_7_port, b => 
                           load_n_store_we_i, outb => n1013);
   U1349 : nand4 port map( a => n520, b => n1014, c => n1015, d => n1016, outb 
                           => n1012);
   U1350 : nor3 port map( a => n1017, b => n1018, c => n1019, outb => n1016);
   U1351 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_5_7_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_1_block_ram_r_3_7_port, d => 
                           n528, outb => n1019);
   U1352 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_7_7_port, b
                           => n529, outb => n1018);
   U1353 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_1_7_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_1_block_ram_r_0_7_port, d => 
                           n531, outb => n1017);
   U1354 : aoi22 port map( a => n532, b => n945, c => n534, d => n959, outb => 
                           n1015);
   U1355 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_2_7_port, 
                           outb => n959);
   U1356 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_4_7_port, 
                           outb => n945);
   U1357 : nand2 port map( a => n536, b => n931, outb => n1014);
   U1358 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_6_7_port, 
                           outb => n931);
   U1359 : nand4 port map( a => n538, b => n1020, c => n1021, d => n1022, outb 
                           => n1011);
   U1360 : nor3 port map( a => n1023, b => n1024, c => n1025, outb => n1022);
   U1361 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_13_7_port,
                           b => n527, c => 
                           load_n_store_RGB_Array_1_block_ram_r_11_7_port, d =>
                           n528, outb => n1025);
   U1362 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_15_7_port, 
                           b => n529, outb => n1024);
   U1363 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_9_7_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_1_block_ram_r_8_7_port, d => 
                           n531, outb => n1023);
   U1364 : aoi22 port map( a => n532, b => n887, c => n534, d => n901, outb => 
                           n1021);
   U1365 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_10_7_port,
                           outb => n901);
   U1366 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_12_7_port,
                           outb => n887);
   U1367 : nand2 port map( a => n536, b => n845, outb => n1020);
   U1368 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_14_7_port,
                           outb => n845);
   U1369 : nand3 port map( a => n1026, b => n1027, c => n1028, outb => n2035);
   U1370 : nand2 port map( a => load_n_store_lazy_in_1_6_port, b => 
                           load_n_store_we_i, outb => n1028);
   U1371 : nand4 port map( a => n520, b => n1029, c => n1030, d => n1031, outb 
                           => n1027);
   U1372 : nor3 port map( a => n1032, b => n1033, c => n1034, outb => n1031);
   U1373 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_5_6_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_1_block_ram_r_3_6_port, d => 
                           n528, outb => n1034);
   U1374 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_7_6_port, b
                           => n529, outb => n1033);
   U1375 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_1_6_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_1_block_ram_r_0_6_port, d => 
                           n531, outb => n1032);
   U1376 : aoi22 port map( a => n532, b => n946, c => n534, d => n960, outb => 
                           n1030);
   U1377 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_2_6_port, 
                           outb => n960);
   U1378 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_4_6_port, 
                           outb => n946);
   U1379 : nand2 port map( a => n536, b => n932, outb => n1029);
   U1380 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_6_6_port, 
                           outb => n932);
   U1381 : nand4 port map( a => n538, b => n1035, c => n1036, d => n1037, outb 
                           => n1026);
   U1382 : nor3 port map( a => n1038, b => n1039, c => n1040, outb => n1037);
   U1383 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_13_6_port,
                           b => n527, c => 
                           load_n_store_RGB_Array_1_block_ram_r_11_6_port, d =>
                           n528, outb => n1040);
   U1384 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_15_6_port, 
                           b => n529, outb => n1039);
   U1385 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_9_6_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_1_block_ram_r_8_6_port, d => 
                           n531, outb => n1038);
   U1386 : aoi22 port map( a => n532, b => n888, c => n534, d => n902, outb => 
                           n1036);
   U1387 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_10_6_port,
                           outb => n902);
   U1388 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_12_6_port,
                           outb => n888);
   U1389 : nand2 port map( a => n536, b => n847, outb => n1035);
   U1390 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_14_6_port,
                           outb => n847);
   U1391 : nand3 port map( a => n1041, b => n1042, c => n1043, outb => n2034);
   U1392 : nand2 port map( a => load_n_store_lazy_in_1_5_port, b => 
                           load_n_store_we_i, outb => n1043);
   U1393 : nand4 port map( a => n520, b => n1044, c => n1045, d => n1046, outb 
                           => n1042);
   U1394 : nor3 port map( a => n1047, b => n1048, c => n1049, outb => n1046);
   U1395 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_5_5_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_1_block_ram_r_3_5_port, d => 
                           n528, outb => n1049);
   U1396 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_7_5_port, b
                           => n529, outb => n1048);
   U1397 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_1_5_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_1_block_ram_r_0_5_port, d => 
                           n531, outb => n1047);
   U1398 : aoi22 port map( a => n532, b => n947, c => n534, d => n961, outb => 
                           n1045);
   U1399 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_2_5_port, 
                           outb => n961);
   U1400 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_4_5_port, 
                           outb => n947);
   U1401 : nand2 port map( a => n536, b => n933, outb => n1044);
   U1402 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_6_5_port, 
                           outb => n933);
   U1403 : nand4 port map( a => n538, b => n1050, c => n1051, d => n1052, outb 
                           => n1041);
   U1404 : nor3 port map( a => n1053, b => n1054, c => n1055, outb => n1052);
   U1405 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_13_5_port,
                           b => n527, c => 
                           load_n_store_RGB_Array_1_block_ram_r_11_5_port, d =>
                           n528, outb => n1055);
   U1406 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_15_5_port, 
                           b => n529, outb => n1054);
   U1407 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_9_5_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_1_block_ram_r_8_5_port, d => 
                           n531, outb => n1053);
   U1408 : aoi22 port map( a => n532, b => n889, c => n534, d => n903, outb => 
                           n1051);
   U1409 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_10_5_port,
                           outb => n903);
   U1410 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_12_5_port,
                           outb => n889);
   U1411 : nand2 port map( a => n536, b => n849, outb => n1050);
   U1412 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_14_5_port,
                           outb => n849);
   U1413 : nand3 port map( a => n1056, b => n1057, c => n1058, outb => n2033);
   U1414 : nand2 port map( a => load_n_store_lazy_in_1_4_port, b => 
                           load_n_store_we_i, outb => n1058);
   U1415 : nand4 port map( a => n520, b => n1059, c => n1060, d => n1061, outb 
                           => n1057);
   U1416 : nor3 port map( a => n1062, b => n1063, c => n1064, outb => n1061);
   U1417 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_5_4_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_1_block_ram_r_3_4_port, d => 
                           n528, outb => n1064);
   U1418 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_7_4_port, b
                           => n529, outb => n1063);
   U1419 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_1_4_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_1_block_ram_r_0_4_port, d => 
                           n531, outb => n1062);
   U1420 : aoi22 port map( a => n532, b => n948, c => n534, d => n962, outb => 
                           n1060);
   U1421 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_2_4_port, 
                           outb => n962);
   U1422 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_4_4_port, 
                           outb => n948);
   U1423 : nand2 port map( a => n536, b => n934, outb => n1059);
   U1424 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_6_4_port, 
                           outb => n934);
   U1425 : nand4 port map( a => n538, b => n1065, c => n1066, d => n1067, outb 
                           => n1056);
   U1426 : nor3 port map( a => n1068, b => n1069, c => n1070, outb => n1067);
   U1427 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_13_4_port,
                           b => n527, c => 
                           load_n_store_RGB_Array_1_block_ram_r_11_4_port, d =>
                           n528, outb => n1070);
   U1428 : nor2 port map( a => load_n_store_RGB_Array_1_block_ram_r_15_4_port, 
                           b => n529, outb => n1069);
   U1429 : oai22 port map( a => load_n_store_RGB_Array_1_block_ram_r_9_4_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_1_block_ram_r_8_4_port, d => 
                           n531, outb => n1068);
   U1430 : aoi22 port map( a => n532, b => n890, c => n534, d => n904, outb => 
                           n1066);
   U1431 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_10_4_port,
                           outb => n904);
   U1432 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_12_4_port,
                           outb => n890);
   U1433 : nand2 port map( a => n536, b => n872, outb => n1065);
   U1434 : inv port map( inb => load_n_store_RGB_Array_1_block_ram_r_14_4_port,
                           outb => n872);
   U1435 : nand3 port map( a => n1071, b => n1072, c => n1073, outb => 
                           load_n_store_RGB_Array_0_n82);
   U1436 : nand2 port map( a => load_n_store_lazy_in_0_3_port, b => 
                           load_n_store_we_i, outb => n1073);
   U1437 : nand4 port map( a => n520, b => n1074, c => n1075, d => n1076, outb 
                           => n1072);
   U1438 : nor3 port map( a => n1077, b => n1078, c => n1079, outb => n1076);
   U1439 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_5_3_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_0_block_ram_r_3_3_port, d => 
                           n528, outb => n1079);
   U1440 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_7_3_port, b
                           => n529, outb => n1078);
   U1441 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_1_3_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_0_block_ram_r_0_3_port, d => 
                           n531, outb => n1077);
   U1442 : aoi22 port map( a => n532, b => n1080, c => n534, d => n1081, outb 
                           => n1075);
   U1443 : nand2 port map( a => n536, b => n1082, outb => n1074);
   U1444 : nand4 port map( a => n538, b => n1083, c => n1084, d => n1085, outb 
                           => n1071);
   U1445 : nor3 port map( a => n1086, b => n1087, c => n1088, outb => n1085);
   U1446 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_13_3_port,
                           b => n527, c => 
                           load_n_store_RGB_Array_0_block_ram_r_11_3_port, d =>
                           n528, outb => n1088);
   U1447 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_15_3_port, 
                           b => n529, outb => n1087);
   U1448 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_9_3_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_0_block_ram_r_8_3_port, d => 
                           n531, outb => n1086);
   U1449 : aoi22 port map( a => n532, b => n1089, c => n534, d => n1090, outb 
                           => n1084);
   U1450 : nand2 port map( a => n536, b => n1091, outb => n1083);
   U1451 : inv port map( inb => n1092, outb => load_n_store_RGB_Array_0_n600);
   U1452 : aoi22 port map( a => load_n_store_lazy_in_0_7_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_0_block_ram_r_15_7_port, outb
                           => n1092);
   U1453 : inv port map( inb => n1093, outb => load_n_store_RGB_Array_0_n599);
   U1454 : aoi22 port map( a => load_n_store_lazy_in_0_6_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_0_block_ram_r_15_6_port, outb
                           => n1093);
   U1455 : inv port map( inb => n1094, outb => load_n_store_RGB_Array_0_n598);
   U1456 : aoi22 port map( a => load_n_store_lazy_in_0_5_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_0_block_ram_r_15_5_port, outb
                           => n1094);
   U1457 : inv port map( inb => n1095, outb => load_n_store_RGB_Array_0_n597);
   U1458 : aoi22 port map( a => load_n_store_lazy_in_0_4_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_0_block_ram_r_15_4_port, outb
                           => n1095);
   U1459 : inv port map( inb => n1096, outb => load_n_store_RGB_Array_0_n596);
   U1460 : aoi22 port map( a => load_n_store_lazy_in_0_3_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_0_block_ram_r_15_3_port, outb
                           => n1096);
   U1461 : inv port map( inb => n1097, outb => load_n_store_RGB_Array_0_n595);
   U1462 : aoi22 port map( a => load_n_store_lazy_in_0_2_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_0_block_ram_r_15_2_port, outb
                           => n1097);
   U1463 : inv port map( inb => n1098, outb => load_n_store_RGB_Array_0_n594);
   U1464 : aoi22 port map( a => load_n_store_lazy_in_0_1_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_0_block_ram_r_15_1_port, outb
                           => n1098);
   U1465 : inv port map( inb => n1099, outb => load_n_store_RGB_Array_0_n593);
   U1466 : aoi22 port map( a => load_n_store_lazy_in_0_0_port, b => n549, c => 
                           n550, d => 
                           load_n_store_RGB_Array_0_block_ram_r_15_0_port, outb
                           => n1099);
   U1467 : inv port map( inb => n550, outb => n549);
   U1468 : nand2 port map( a => n1100, b => n1101, outb => n550);
   U1469 : oai22 port map( a => n1102, b => n559, c => n560, d => n1103, outb 
                           => load_n_store_RGB_Array_0_n592);
   U1470 : oai22 port map( a => n1104, b => n559, c => n560, d => n1105, outb 
                           => load_n_store_RGB_Array_0_n591);
   U1471 : oai22 port map( a => n1106, b => n559, c => n560, d => n1107, outb 
                           => load_n_store_RGB_Array_0_n590);
   U1472 : nand3 port map( a => n1108, b => n1109, c => n1110, outb => 
                           load_n_store_RGB_Array_0_n59);
   U1473 : nand2 port map( a => load_n_store_lazy_in_0_2_port, b => 
                           load_n_store_we_i, outb => n1110);
   U1474 : nand4 port map( a => n520, b => n1111, c => n1112, d => n1113, outb 
                           => n1109);
   U1475 : nor3 port map( a => n1114, b => n1115, c => n1116, outb => n1113);
   U1476 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_5_2_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_0_block_ram_r_3_2_port, d => 
                           n528, outb => n1116);
   U1477 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_7_2_port, b
                           => n529, outb => n1115);
   U1478 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_1_2_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_0_block_ram_r_0_2_port, d => 
                           n531, outb => n1114);
   U1479 : aoi22 port map( a => n532, b => n1117, c => n534, d => n1118, outb 
                           => n1112);
   U1480 : nand2 port map( a => n536, b => n1119, outb => n1111);
   U1481 : nand4 port map( a => n538, b => n1120, c => n1121, d => n1122, outb 
                           => n1108);
   U1482 : nor3 port map( a => n1123, b => n1124, c => n1125, outb => n1122);
   U1483 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_13_2_port,
                           b => n527, c => 
                           load_n_store_RGB_Array_0_block_ram_r_11_2_port, d =>
                           n528, outb => n1125);
   U1484 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_15_2_port, 
                           b => n529, outb => n1124);
   U1485 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_9_2_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_0_block_ram_r_8_2_port, d => 
                           n531, outb => n1123);
   U1486 : aoi22 port map( a => n532, b => n1126, c => n534, d => n1127, outb 
                           => n1121);
   U1487 : nand2 port map( a => n536, b => n1128, outb => n1120);
   U1488 : oai22 port map( a => n1129, b => n559, c => n560, d => n1130, outb 
                           => load_n_store_RGB_Array_0_n589);
   U1489 : oai22 port map( a => n1131, b => n559, c => n560, d => n1091, outb 
                           => load_n_store_RGB_Array_0_n588);
   U1490 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_14_3_port,
                           outb => n1091);
   U1491 : oai22 port map( a => n1132, b => n559, c => n560, d => n1128, outb 
                           => load_n_store_RGB_Array_0_n587);
   U1492 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_14_2_port,
                           outb => n1128);
   U1493 : oai22 port map( a => n1133, b => n559, c => n560, d => n1134, outb 
                           => load_n_store_RGB_Array_0_n586);
   U1494 : oai22 port map( a => n1135, b => n559, c => n560, d => n1136, outb 
                           => load_n_store_RGB_Array_0_n585);
   U1495 : inv port map( inb => n559, outb => n560);
   U1496 : nand2 port map( a => n1100, b => n536, outb => n559);
   U1497 : inv port map( inb => n1137, outb => load_n_store_RGB_Array_0_n584);
   U1498 : aoi22 port map( a => load_n_store_lazy_in_0_7_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_0_block_ram_r_13_7_port, outb
                           => n1137);
   U1499 : inv port map( inb => n1138, outb => load_n_store_RGB_Array_0_n583);
   U1500 : aoi22 port map( a => load_n_store_lazy_in_0_6_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_0_block_ram_r_13_6_port, outb
                           => n1138);
   U1501 : inv port map( inb => n1139, outb => load_n_store_RGB_Array_0_n582);
   U1502 : aoi22 port map( a => load_n_store_lazy_in_0_5_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_0_block_ram_r_13_5_port, outb
                           => n1139);
   U1503 : inv port map( inb => n1140, outb => load_n_store_RGB_Array_0_n581);
   U1504 : aoi22 port map( a => load_n_store_lazy_in_0_4_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_0_block_ram_r_13_4_port, outb
                           => n1140);
   U1505 : inv port map( inb => n1141, outb => load_n_store_RGB_Array_0_n580);
   U1506 : aoi22 port map( a => load_n_store_lazy_in_0_3_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_0_block_ram_r_13_3_port, outb
                           => n1141);
   U1507 : inv port map( inb => n1142, outb => load_n_store_RGB_Array_0_n579);
   U1508 : aoi22 port map( a => load_n_store_lazy_in_0_2_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_0_block_ram_r_13_2_port, outb
                           => n1142);
   U1509 : inv port map( inb => n1143, outb => load_n_store_RGB_Array_0_n578);
   U1510 : aoi22 port map( a => load_n_store_lazy_in_0_1_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_0_block_ram_r_13_1_port, outb
                           => n1143);
   U1511 : inv port map( inb => n1144, outb => load_n_store_RGB_Array_0_n577);
   U1512 : aoi22 port map( a => load_n_store_lazy_in_0_0_port, b => n596, c => 
                           n597, d => 
                           load_n_store_RGB_Array_0_block_ram_r_13_0_port, outb
                           => n1144);
   U1513 : inv port map( inb => n597, outb => n596);
   U1514 : nand2 port map( a => n1100, b => n1145, outb => n597);
   U1515 : oai22 port map( a => n1102, b => n605, c => n606, d => n1146, outb 
                           => load_n_store_RGB_Array_0_n576);
   U1516 : oai22 port map( a => n1104, b => n605, c => n606, d => n1147, outb 
                           => load_n_store_RGB_Array_0_n575);
   U1517 : oai22 port map( a => n1106, b => n605, c => n606, d => n1148, outb 
                           => load_n_store_RGB_Array_0_n574);
   U1518 : oai22 port map( a => n1129, b => n605, c => n606, d => n1149, outb 
                           => load_n_store_RGB_Array_0_n573);
   U1519 : oai22 port map( a => n1131, b => n605, c => n606, d => n1089, outb 
                           => load_n_store_RGB_Array_0_n572);
   U1520 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_12_3_port,
                           outb => n1089);
   U1521 : oai22 port map( a => n1132, b => n605, c => n606, d => n1126, outb 
                           => load_n_store_RGB_Array_0_n571);
   U1522 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_12_2_port,
                           outb => n1126);
   U1523 : oai22 port map( a => n1133, b => n605, c => n606, d => n1150, outb 
                           => load_n_store_RGB_Array_0_n570);
   U1524 : oai22 port map( a => n1135, b => n605, c => n606, d => n1151, outb 
                           => load_n_store_RGB_Array_0_n569);
   U1525 : inv port map( inb => n605, outb => n606);
   U1526 : nand2 port map( a => n1100, b => n532, outb => n605);
   U1527 : inv port map( inb => n1152, outb => load_n_store_RGB_Array_0_n568);
   U1528 : aoi22 port map( a => load_n_store_lazy_in_0_7_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_0_block_ram_r_11_7_port, outb
                           => n1152);
   U1529 : inv port map( inb => n1153, outb => load_n_store_RGB_Array_0_n567);
   U1530 : aoi22 port map( a => load_n_store_lazy_in_0_6_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_0_block_ram_r_11_6_port, outb
                           => n1153);
   U1531 : inv port map( inb => n1154, outb => load_n_store_RGB_Array_0_n566);
   U1532 : aoi22 port map( a => load_n_store_lazy_in_0_5_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_0_block_ram_r_11_5_port, outb
                           => n1154);
   U1533 : inv port map( inb => n1155, outb => load_n_store_RGB_Array_0_n565);
   U1534 : aoi22 port map( a => load_n_store_lazy_in_0_4_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_0_block_ram_r_11_4_port, outb
                           => n1155);
   U1535 : inv port map( inb => n1156, outb => load_n_store_RGB_Array_0_n564);
   U1536 : aoi22 port map( a => load_n_store_lazy_in_0_3_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_0_block_ram_r_11_3_port, outb
                           => n1156);
   U1537 : inv port map( inb => n1157, outb => load_n_store_RGB_Array_0_n563);
   U1538 : aoi22 port map( a => load_n_store_lazy_in_0_2_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_0_block_ram_r_11_2_port, outb
                           => n1157);
   U1539 : inv port map( inb => n1158, outb => load_n_store_RGB_Array_0_n562);
   U1540 : aoi22 port map( a => load_n_store_lazy_in_0_1_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_0_block_ram_r_11_1_port, outb
                           => n1158);
   U1541 : inv port map( inb => n1159, outb => load_n_store_RGB_Array_0_n561);
   U1542 : aoi22 port map( a => load_n_store_lazy_in_0_0_port, b => n614, c => 
                           n615, d => 
                           load_n_store_RGB_Array_0_block_ram_r_11_0_port, outb
                           => n1159);
   U1543 : inv port map( inb => n615, outb => n614);
   U1544 : nand2 port map( a => n1100, b => n1160, outb => n615);
   U1545 : oai22 port map( a => n1102, b => n623, c => n624, d => n1161, outb 
                           => load_n_store_RGB_Array_0_n560);
   U1546 : oai22 port map( a => n1104, b => n623, c => n624, d => n1162, outb 
                           => load_n_store_RGB_Array_0_n559);
   U1547 : oai22 port map( a => n1106, b => n623, c => n624, d => n1163, outb 
                           => load_n_store_RGB_Array_0_n558);
   U1548 : oai22 port map( a => n1129, b => n623, c => n624, d => n1164, outb 
                           => load_n_store_RGB_Array_0_n557);
   U1549 : oai22 port map( a => n1131, b => n623, c => n624, d => n1090, outb 
                           => load_n_store_RGB_Array_0_n556);
   U1550 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_10_3_port,
                           outb => n1090);
   U1551 : oai22 port map( a => n1132, b => n623, c => n624, d => n1127, outb 
                           => load_n_store_RGB_Array_0_n555);
   U1552 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_10_2_port,
                           outb => n1127);
   U1553 : oai22 port map( a => n1133, b => n623, c => n624, d => n1165, outb 
                           => load_n_store_RGB_Array_0_n554);
   U1554 : oai22 port map( a => n1135, b => n623, c => n624, d => n1166, outb 
                           => load_n_store_RGB_Array_0_n553);
   U1555 : inv port map( inb => n623, outb => n624);
   U1556 : nand2 port map( a => n1100, b => n534, outb => n623);
   U1557 : inv port map( inb => n1167, outb => load_n_store_RGB_Array_0_n552);
   U1558 : aoi22 port map( a => load_n_store_lazy_in_0_7_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_0_block_ram_r_9_7_port, outb 
                           => n1167);
   U1559 : inv port map( inb => n1168, outb => load_n_store_RGB_Array_0_n551);
   U1560 : aoi22 port map( a => load_n_store_lazy_in_0_6_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_0_block_ram_r_9_6_port, outb 
                           => n1168);
   U1561 : inv port map( inb => n1169, outb => load_n_store_RGB_Array_0_n550);
   U1562 : aoi22 port map( a => load_n_store_lazy_in_0_5_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_0_block_ram_r_9_5_port, outb 
                           => n1169);
   U1563 : inv port map( inb => n1170, outb => load_n_store_RGB_Array_0_n549);
   U1564 : aoi22 port map( a => load_n_store_lazy_in_0_4_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_0_block_ram_r_9_4_port, outb 
                           => n1170);
   U1565 : inv port map( inb => n1171, outb => load_n_store_RGB_Array_0_n548);
   U1566 : aoi22 port map( a => load_n_store_lazy_in_0_3_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_0_block_ram_r_9_3_port, outb 
                           => n1171);
   U1567 : inv port map( inb => n1172, outb => load_n_store_RGB_Array_0_n547);
   U1568 : aoi22 port map( a => load_n_store_lazy_in_0_2_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_0_block_ram_r_9_2_port, outb 
                           => n1172);
   U1569 : inv port map( inb => n1173, outb => load_n_store_RGB_Array_0_n546);
   U1570 : aoi22 port map( a => load_n_store_lazy_in_0_1_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_0_block_ram_r_9_1_port, outb 
                           => n1173);
   U1571 : inv port map( inb => n1174, outb => load_n_store_RGB_Array_0_n545);
   U1572 : aoi22 port map( a => load_n_store_lazy_in_0_0_port, b => n632, c => 
                           n633, d => 
                           load_n_store_RGB_Array_0_block_ram_r_9_0_port, outb 
                           => n1174);
   U1573 : inv port map( inb => n633, outb => n632);
   U1574 : nand2 port map( a => n1100, b => n1175, outb => n633);
   U1575 : inv port map( inb => n1176, outb => load_n_store_RGB_Array_0_n544);
   U1576 : aoi22 port map( a => load_n_store_lazy_in_0_7_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_0_block_ram_r_8_7_port, outb 
                           => n1176);
   U1577 : inv port map( inb => n1177, outb => load_n_store_RGB_Array_0_n543);
   U1578 : aoi22 port map( a => load_n_store_lazy_in_0_6_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_0_block_ram_r_8_6_port, outb 
                           => n1177);
   U1579 : inv port map( inb => n1178, outb => load_n_store_RGB_Array_0_n542);
   U1580 : aoi22 port map( a => load_n_store_lazy_in_0_5_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_0_block_ram_r_8_5_port, outb 
                           => n1178);
   U1581 : inv port map( inb => n1179, outb => load_n_store_RGB_Array_0_n541);
   U1582 : aoi22 port map( a => load_n_store_lazy_in_0_4_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_0_block_ram_r_8_4_port, outb 
                           => n1179);
   U1583 : inv port map( inb => n1180, outb => load_n_store_RGB_Array_0_n540);
   U1584 : aoi22 port map( a => load_n_store_lazy_in_0_3_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_0_block_ram_r_8_3_port, outb 
                           => n1180);
   U1585 : inv port map( inb => n1181, outb => load_n_store_RGB_Array_0_n539);
   U1586 : aoi22 port map( a => load_n_store_lazy_in_0_2_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_0_block_ram_r_8_2_port, outb 
                           => n1181);
   U1587 : inv port map( inb => n1182, outb => load_n_store_RGB_Array_0_n538);
   U1588 : aoi22 port map( a => load_n_store_lazy_in_0_1_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_0_block_ram_r_8_1_port, outb 
                           => n1182);
   U1589 : inv port map( inb => n1183, outb => load_n_store_RGB_Array_0_n537);
   U1590 : aoi22 port map( a => load_n_store_lazy_in_0_0_port, b => n642, c => 
                           n643, d => 
                           load_n_store_RGB_Array_0_block_ram_r_8_0_port, outb 
                           => n1183);
   U1591 : inv port map( inb => n643, outb => n642);
   U1592 : nand2 port map( a => n1100, b => n1184, outb => n643);
   U1593 : nor2 port map( a => n136, b => n46, outb => n1100);
   U1594 : inv port map( inb => n1185, outb => load_n_store_RGB_Array_0_n536);
   U1595 : aoi22 port map( a => load_n_store_lazy_in_0_7_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_0_block_ram_r_7_7_port, outb 
                           => n1185);
   U1596 : inv port map( inb => n1186, outb => load_n_store_RGB_Array_0_n535);
   U1597 : aoi22 port map( a => load_n_store_lazy_in_0_6_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_0_block_ram_r_7_6_port, outb 
                           => n1186);
   U1598 : inv port map( inb => n1187, outb => load_n_store_RGB_Array_0_n534);
   U1599 : aoi22 port map( a => load_n_store_lazy_in_0_5_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_0_block_ram_r_7_5_port, outb 
                           => n1187);
   U1600 : inv port map( inb => n1188, outb => load_n_store_RGB_Array_0_n533);
   U1601 : aoi22 port map( a => load_n_store_lazy_in_0_4_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_0_block_ram_r_7_4_port, outb 
                           => n1188);
   U1602 : inv port map( inb => n1189, outb => load_n_store_RGB_Array_0_n532);
   U1603 : aoi22 port map( a => load_n_store_lazy_in_0_3_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_0_block_ram_r_7_3_port, outb 
                           => n1189);
   U1604 : inv port map( inb => n1190, outb => load_n_store_RGB_Array_0_n531);
   U1605 : aoi22 port map( a => load_n_store_lazy_in_0_2_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_0_block_ram_r_7_2_port, outb 
                           => n1190);
   U1606 : inv port map( inb => n1191, outb => load_n_store_RGB_Array_0_n530);
   U1607 : aoi22 port map( a => load_n_store_lazy_in_0_1_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_0_block_ram_r_7_1_port, outb 
                           => n1191);
   U1608 : inv port map( inb => n1192, outb => load_n_store_RGB_Array_0_n529);
   U1609 : aoi22 port map( a => load_n_store_lazy_in_0_0_port, b => n652, c => 
                           n653, d => 
                           load_n_store_RGB_Array_0_block_ram_r_7_0_port, outb 
                           => n1192);
   U1610 : inv port map( inb => n653, outb => n652);
   U1611 : nand2 port map( a => n1193, b => n1101, outb => n653);
   U1612 : oai22 port map( a => n1102, b => n661, c => n662, d => n1194, outb 
                           => load_n_store_RGB_Array_0_n528);
   U1613 : oai22 port map( a => n1104, b => n661, c => n662, d => n1195, outb 
                           => load_n_store_RGB_Array_0_n527);
   U1614 : oai22 port map( a => n1106, b => n661, c => n662, d => n1196, outb 
                           => load_n_store_RGB_Array_0_n526);
   U1615 : oai22 port map( a => n1129, b => n661, c => n662, d => n1197, outb 
                           => load_n_store_RGB_Array_0_n525);
   U1616 : oai22 port map( a => n1131, b => n661, c => n662, d => n1082, outb 
                           => load_n_store_RGB_Array_0_n524);
   U1617 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_6_3_port, 
                           outb => n1082);
   U1618 : oai22 port map( a => n1132, b => n661, c => n662, d => n1119, outb 
                           => load_n_store_RGB_Array_0_n523);
   U1619 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_6_2_port, 
                           outb => n1119);
   U1620 : oai22 port map( a => n1133, b => n661, c => n662, d => n1198, outb 
                           => load_n_store_RGB_Array_0_n522);
   U1621 : oai22 port map( a => n1135, b => n661, c => n662, d => n1199, outb 
                           => load_n_store_RGB_Array_0_n521);
   U1622 : inv port map( inb => n661, outb => n662);
   U1623 : nand2 port map( a => n1193, b => n536, outb => n661);
   U1624 : inv port map( inb => n1200, outb => load_n_store_RGB_Array_0_n520);
   U1625 : aoi22 port map( a => load_n_store_lazy_in_0_7_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_0_block_ram_r_5_7_port, outb 
                           => n1200);
   U1626 : inv port map( inb => n1201, outb => load_n_store_RGB_Array_0_n519);
   U1627 : aoi22 port map( a => load_n_store_lazy_in_0_6_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_0_block_ram_r_5_6_port, outb 
                           => n1201);
   U1628 : inv port map( inb => n1202, outb => load_n_store_RGB_Array_0_n518);
   U1629 : aoi22 port map( a => load_n_store_lazy_in_0_5_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_0_block_ram_r_5_5_port, outb 
                           => n1202);
   U1630 : inv port map( inb => n1203, outb => load_n_store_RGB_Array_0_n517);
   U1631 : aoi22 port map( a => load_n_store_lazy_in_0_4_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_0_block_ram_r_5_4_port, outb 
                           => n1203);
   U1632 : inv port map( inb => n1204, outb => load_n_store_RGB_Array_0_n516);
   U1633 : aoi22 port map( a => load_n_store_lazy_in_0_3_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_0_block_ram_r_5_3_port, outb 
                           => n1204);
   U1634 : inv port map( inb => n1205, outb => load_n_store_RGB_Array_0_n515);
   U1635 : aoi22 port map( a => load_n_store_lazy_in_0_2_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_0_block_ram_r_5_2_port, outb 
                           => n1205);
   U1636 : inv port map( inb => n1206, outb => load_n_store_RGB_Array_0_n514);
   U1637 : aoi22 port map( a => load_n_store_lazy_in_0_1_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_0_block_ram_r_5_1_port, outb 
                           => n1206);
   U1638 : inv port map( inb => n1207, outb => load_n_store_RGB_Array_0_n513);
   U1639 : aoi22 port map( a => load_n_store_lazy_in_0_0_port, b => n670, c => 
                           n671, d => 
                           load_n_store_RGB_Array_0_block_ram_r_5_0_port, outb 
                           => n1207);
   U1640 : inv port map( inb => n671, outb => n670);
   U1641 : nand2 port map( a => n1193, b => n1145, outb => n671);
   U1642 : oai22 port map( a => n1102, b => n679, c => n680, d => n1208, outb 
                           => load_n_store_RGB_Array_0_n512);
   U1643 : oai22 port map( a => n1104, b => n679, c => n680, d => n1209, outb 
                           => load_n_store_RGB_Array_0_n511);
   U1644 : oai22 port map( a => n1106, b => n679, c => n680, d => n1210, outb 
                           => load_n_store_RGB_Array_0_n510);
   U1645 : oai22 port map( a => n1129, b => n679, c => n680, d => n1211, outb 
                           => load_n_store_RGB_Array_0_n509);
   U1646 : oai22 port map( a => n1131, b => n679, c => n680, d => n1080, outb 
                           => load_n_store_RGB_Array_0_n508);
   U1647 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_4_3_port, 
                           outb => n1080);
   U1648 : oai22 port map( a => n1132, b => n679, c => n680, d => n1117, outb 
                           => load_n_store_RGB_Array_0_n507);
   U1649 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_4_2_port, 
                           outb => n1117);
   U1650 : oai22 port map( a => n1133, b => n679, c => n680, d => n1212, outb 
                           => load_n_store_RGB_Array_0_n506);
   U1651 : oai22 port map( a => n1135, b => n679, c => n680, d => n1213, outb 
                           => load_n_store_RGB_Array_0_n505);
   U1652 : inv port map( inb => n679, outb => n680);
   U1653 : nand2 port map( a => n1193, b => n532, outb => n679);
   U1654 : inv port map( inb => n1214, outb => load_n_store_RGB_Array_0_n504);
   U1655 : aoi22 port map( a => load_n_store_lazy_in_0_7_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_0_block_ram_r_3_7_port, outb 
                           => n1214);
   U1656 : inv port map( inb => n1215, outb => load_n_store_RGB_Array_0_n503);
   U1657 : aoi22 port map( a => load_n_store_lazy_in_0_6_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_0_block_ram_r_3_6_port, outb 
                           => n1215);
   U1658 : inv port map( inb => n1216, outb => load_n_store_RGB_Array_0_n502);
   U1659 : aoi22 port map( a => load_n_store_lazy_in_0_5_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_0_block_ram_r_3_5_port, outb 
                           => n1216);
   U1660 : inv port map( inb => n1217, outb => load_n_store_RGB_Array_0_n501);
   U1661 : aoi22 port map( a => load_n_store_lazy_in_0_4_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_0_block_ram_r_3_4_port, outb 
                           => n1217);
   U1662 : inv port map( inb => n1218, outb => load_n_store_RGB_Array_0_n500);
   U1663 : aoi22 port map( a => load_n_store_lazy_in_0_3_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_0_block_ram_r_3_3_port, outb 
                           => n1218);
   U1664 : inv port map( inb => n1219, outb => load_n_store_RGB_Array_0_n499);
   U1665 : aoi22 port map( a => load_n_store_lazy_in_0_2_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_0_block_ram_r_3_2_port, outb 
                           => n1219);
   U1666 : inv port map( inb => n1220, outb => load_n_store_RGB_Array_0_n498);
   U1667 : aoi22 port map( a => load_n_store_lazy_in_0_1_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_0_block_ram_r_3_1_port, outb 
                           => n1220);
   U1668 : inv port map( inb => n1221, outb => load_n_store_RGB_Array_0_n497);
   U1669 : aoi22 port map( a => load_n_store_lazy_in_0_0_port, b => n688, c => 
                           n689, d => 
                           load_n_store_RGB_Array_0_block_ram_r_3_0_port, outb 
                           => n1221);
   U1670 : inv port map( inb => n689, outb => n688);
   U1671 : nand2 port map( a => n1193, b => n1160, outb => n689);
   U1672 : oai22 port map( a => n1102, b => n697, c => n698, d => n1222, outb 
                           => load_n_store_RGB_Array_0_n496);
   U1673 : inv port map( inb => load_n_store_lazy_in_0_7_port, outb => n1102);
   U1674 : oai22 port map( a => n1104, b => n697, c => n698, d => n1223, outb 
                           => load_n_store_RGB_Array_0_n495);
   U1675 : inv port map( inb => load_n_store_lazy_in_0_6_port, outb => n1104);
   U1676 : oai22 port map( a => n1106, b => n697, c => n698, d => n1224, outb 
                           => load_n_store_RGB_Array_0_n494);
   U1677 : inv port map( inb => load_n_store_lazy_in_0_5_port, outb => n1106);
   U1678 : oai22 port map( a => n1129, b => n697, c => n698, d => n1225, outb 
                           => load_n_store_RGB_Array_0_n493);
   U1679 : inv port map( inb => load_n_store_lazy_in_0_4_port, outb => n1129);
   U1680 : oai22 port map( a => n1131, b => n697, c => n698, d => n1081, outb 
                           => load_n_store_RGB_Array_0_n492);
   U1681 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_2_3_port, 
                           outb => n1081);
   U1682 : inv port map( inb => load_n_store_lazy_in_0_3_port, outb => n1131);
   U1683 : oai22 port map( a => n1132, b => n697, c => n698, d => n1118, outb 
                           => load_n_store_RGB_Array_0_n491);
   U1684 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_2_2_port, 
                           outb => n1118);
   U1685 : inv port map( inb => load_n_store_lazy_in_0_2_port, outb => n1132);
   U1686 : oai22 port map( a => n1133, b => n697, c => n698, d => n1226, outb 
                           => load_n_store_RGB_Array_0_n490);
   U1687 : inv port map( inb => load_n_store_lazy_in_0_1_port, outb => n1133);
   U1688 : oai22 port map( a => n1135, b => n697, c => n698, d => n1227, outb 
                           => load_n_store_RGB_Array_0_n489);
   U1689 : inv port map( inb => n697, outb => n698);
   U1690 : nand2 port map( a => n1193, b => n534, outb => n697);
   U1691 : inv port map( inb => load_n_store_lazy_in_0_0_port, outb => n1135);
   U1692 : inv port map( inb => n1228, outb => load_n_store_RGB_Array_0_n488);
   U1693 : aoi22 port map( a => load_n_store_lazy_in_0_7_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_0_block_ram_r_1_7_port, outb 
                           => n1228);
   U1694 : inv port map( inb => n1229, outb => load_n_store_RGB_Array_0_n487);
   U1695 : aoi22 port map( a => load_n_store_lazy_in_0_6_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_0_block_ram_r_1_6_port, outb 
                           => n1229);
   U1696 : inv port map( inb => n1230, outb => load_n_store_RGB_Array_0_n486);
   U1697 : aoi22 port map( a => load_n_store_lazy_in_0_5_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_0_block_ram_r_1_5_port, outb 
                           => n1230);
   U1698 : inv port map( inb => n1231, outb => load_n_store_RGB_Array_0_n485);
   U1699 : aoi22 port map( a => load_n_store_lazy_in_0_4_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_0_block_ram_r_1_4_port, outb 
                           => n1231);
   U1700 : inv port map( inb => n1232, outb => load_n_store_RGB_Array_0_n484);
   U1701 : aoi22 port map( a => load_n_store_lazy_in_0_3_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_0_block_ram_r_1_3_port, outb 
                           => n1232);
   U1702 : inv port map( inb => n1233, outb => load_n_store_RGB_Array_0_n483);
   U1703 : aoi22 port map( a => load_n_store_lazy_in_0_2_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_0_block_ram_r_1_2_port, outb 
                           => n1233);
   U1704 : inv port map( inb => n1234, outb => load_n_store_RGB_Array_0_n482);
   U1705 : aoi22 port map( a => load_n_store_lazy_in_0_1_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_0_block_ram_r_1_1_port, outb 
                           => n1234);
   U1706 : inv port map( inb => n1235, outb => load_n_store_RGB_Array_0_n481);
   U1707 : aoi22 port map( a => load_n_store_lazy_in_0_0_port, b => n706, c => 
                           n707, d => 
                           load_n_store_RGB_Array_0_block_ram_r_1_0_port, outb 
                           => n1235);
   U1708 : inv port map( inb => n707, outb => n706);
   U1709 : nand2 port map( a => n1193, b => n1175, outb => n707);
   U1710 : inv port map( inb => n1236, outb => load_n_store_RGB_Array_0_n480);
   U1711 : aoi22 port map( a => load_n_store_lazy_in_0_7_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_0_block_ram_r_0_7_port, outb 
                           => n1236);
   U1712 : inv port map( inb => n1237, outb => load_n_store_RGB_Array_0_n479);
   U1713 : aoi22 port map( a => load_n_store_lazy_in_0_6_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_0_block_ram_r_0_6_port, outb 
                           => n1237);
   U1714 : inv port map( inb => n1238, outb => load_n_store_RGB_Array_0_n478);
   U1715 : aoi22 port map( a => load_n_store_lazy_in_0_5_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_0_block_ram_r_0_5_port, outb 
                           => n1238);
   U1716 : inv port map( inb => n1239, outb => load_n_store_RGB_Array_0_n477);
   U1717 : aoi22 port map( a => load_n_store_lazy_in_0_4_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_0_block_ram_r_0_4_port, outb 
                           => n1239);
   U1718 : inv port map( inb => n1240, outb => load_n_store_RGB_Array_0_n476);
   U1719 : aoi22 port map( a => load_n_store_lazy_in_0_3_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_0_block_ram_r_0_3_port, outb 
                           => n1240);
   U1720 : inv port map( inb => n1241, outb => load_n_store_RGB_Array_0_n475);
   U1721 : aoi22 port map( a => load_n_store_lazy_in_0_2_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_0_block_ram_r_0_2_port, outb 
                           => n1241);
   U1722 : inv port map( inb => n1242, outb => load_n_store_RGB_Array_0_n474);
   U1723 : aoi22 port map( a => load_n_store_lazy_in_0_1_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_0_block_ram_r_0_1_port, outb 
                           => n1242);
   U1724 : inv port map( inb => n1243, outb => load_n_store_RGB_Array_0_n473);
   U1725 : aoi22 port map( a => load_n_store_lazy_in_0_0_port, b => n716, c => 
                           n717, d => 
                           load_n_store_RGB_Array_0_block_ram_r_0_0_port, outb 
                           => n1243);
   U1726 : inv port map( inb => n717, outb => n716);
   U1727 : nand2 port map( a => n1193, b => n1184, outb => n717);
   U1728 : nor2 port map( a => n136, b => addr_i_3_port, outb => n1193);
   U1729 : inv port map( inb => load_n_store_we_i, outb => n136);
   U1730 : nand3 port map( a => n1244, b => n1245, c => n1246, outb => 
                           load_n_store_RGB_Array_0_n36);
   U1731 : nand2 port map( a => load_n_store_lazy_in_0_1_port, b => 
                           load_n_store_we_i, outb => n1246);
   U1732 : nand4 port map( a => n520, b => n1247, c => n1248, d => n1249, outb 
                           => n1245);
   U1733 : nor3 port map( a => n1250, b => n1251, c => n1252, outb => n1249);
   U1734 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_5_1_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_0_block_ram_r_3_1_port, d => 
                           n528, outb => n1252);
   U1735 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_7_1_port, b
                           => n529, outb => n1251);
   U1736 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_1_1_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_0_block_ram_r_0_1_port, d => 
                           n531, outb => n1250);
   U1737 : aoi22 port map( a => n532, b => n1212, c => n534, d => n1226, outb 
                           => n1248);
   U1738 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_2_1_port, 
                           outb => n1226);
   U1739 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_4_1_port, 
                           outb => n1212);
   U1740 : nand2 port map( a => n536, b => n1198, outb => n1247);
   U1741 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_6_1_port, 
                           outb => n1198);
   U1742 : nand4 port map( a => n538, b => n1253, c => n1254, d => n1255, outb 
                           => n1244);
   U1743 : nor3 port map( a => n1256, b => n1257, c => n1258, outb => n1255);
   U1744 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_13_1_port,
                           b => n527, c => 
                           load_n_store_RGB_Array_0_block_ram_r_11_1_port, d =>
                           n528, outb => n1258);
   U1745 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_15_1_port, 
                           b => n529, outb => n1257);
   U1746 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_9_1_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_0_block_ram_r_8_1_port, d => 
                           n531, outb => n1256);
   U1747 : aoi22 port map( a => n532, b => n1150, c => n534, d => n1165, outb 
                           => n1254);
   U1748 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_10_1_port,
                           outb => n1165);
   U1749 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_12_1_port,
                           outb => n1150);
   U1750 : nand2 port map( a => n536, b => n1134, outb => n1253);
   U1751 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_14_1_port,
                           outb => n1134);
   U1752 : nand3 port map( a => n1259, b => n1260, c => n1261, outb => 
                           load_n_store_RGB_Array_0_n2);
   U1753 : nand2 port map( a => load_n_store_lazy_in_0_0_port, b => 
                           load_n_store_we_i, outb => n1261);
   U1754 : nand4 port map( a => n520, b => n1262, c => n1263, d => n1264, outb 
                           => n1260);
   U1755 : nor3 port map( a => n1265, b => n1266, c => n1267, outb => n1264);
   U1756 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_5_0_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_0_block_ram_r_3_0_port, d => 
                           n528, outb => n1267);
   U1757 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_7_0_port, b
                           => n529, outb => n1266);
   U1758 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_1_0_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_0_block_ram_r_0_0_port, d => 
                           n531, outb => n1265);
   U1759 : aoi22 port map( a => n532, b => n1213, c => n534, d => n1227, outb 
                           => n1263);
   U1760 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_2_0_port, 
                           outb => n1227);
   U1761 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_4_0_port, 
                           outb => n1213);
   U1762 : nand2 port map( a => n536, b => n1199, outb => n1262);
   U1763 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_6_0_port, 
                           outb => n1199);
   U1764 : nand4 port map( a => n538, b => n1268, c => n1269, d => n1270, outb 
                           => n1259);
   U1765 : nor3 port map( a => n1271, b => n1272, c => n1273, outb => n1270);
   U1766 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_13_0_port,
                           b => n527, c => 
                           load_n_store_RGB_Array_0_block_ram_r_11_0_port, d =>
                           n528, outb => n1273);
   U1767 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_15_0_port, 
                           b => n529, outb => n1272);
   U1768 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_9_0_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_0_block_ram_r_8_0_port, d => 
                           n531, outb => n1271);
   U1769 : aoi22 port map( a => n532, b => n1151, c => n534, d => n1166, outb 
                           => n1269);
   U1770 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_10_0_port,
                           outb => n1166);
   U1771 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_12_0_port,
                           outb => n1151);
   U1772 : nand2 port map( a => n536, b => n1136, outb => n1268);
   U1773 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_14_0_port,
                           outb => n1136);
   U1774 : nand3 port map( a => n1274, b => n1275, c => n1276, outb => 
                           load_n_store_RGB_Array_0_n174);
   U1775 : nand2 port map( a => load_n_store_lazy_in_0_7_port, b => 
                           load_n_store_we_i, outb => n1276);
   U1776 : nand4 port map( a => n520, b => n1277, c => n1278, d => n1279, outb 
                           => n1275);
   U1777 : nor3 port map( a => n1280, b => n1281, c => n1282, outb => n1279);
   U1778 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_5_7_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_0_block_ram_r_3_7_port, d => 
                           n528, outb => n1282);
   U1779 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_7_7_port, b
                           => n529, outb => n1281);
   U1780 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_1_7_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_0_block_ram_r_0_7_port, d => 
                           n531, outb => n1280);
   U1781 : aoi22 port map( a => n532, b => n1208, c => n534, d => n1222, outb 
                           => n1278);
   U1782 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_2_7_port, 
                           outb => n1222);
   U1783 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_4_7_port, 
                           outb => n1208);
   U1784 : nand2 port map( a => n536, b => n1194, outb => n1277);
   U1785 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_6_7_port, 
                           outb => n1194);
   U1786 : nand4 port map( a => n538, b => n1283, c => n1284, d => n1285, outb 
                           => n1274);
   U1787 : nor3 port map( a => n1286, b => n1287, c => n1288, outb => n1285);
   U1788 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_13_7_port,
                           b => n527, c => 
                           load_n_store_RGB_Array_0_block_ram_r_11_7_port, d =>
                           n528, outb => n1288);
   U1789 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_15_7_port, 
                           b => n529, outb => n1287);
   U1790 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_9_7_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_0_block_ram_r_8_7_port, d => 
                           n531, outb => n1286);
   U1791 : aoi22 port map( a => n532, b => n1146, c => n534, d => n1161, outb 
                           => n1284);
   U1792 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_10_7_port,
                           outb => n1161);
   U1793 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_12_7_port,
                           outb => n1146);
   U1794 : nand2 port map( a => n536, b => n1103, outb => n1283);
   U1795 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_14_7_port,
                           outb => n1103);
   U1796 : nand3 port map( a => n1289, b => n1290, c => n1291, outb => 
                           load_n_store_RGB_Array_0_n151);
   U1797 : nand2 port map( a => load_n_store_lazy_in_0_6_port, b => 
                           load_n_store_we_i, outb => n1291);
   U1798 : nand4 port map( a => n520, b => n1292, c => n1293, d => n1294, outb 
                           => n1290);
   U1799 : nor3 port map( a => n1295, b => n1296, c => n1297, outb => n1294);
   U1800 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_5_6_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_0_block_ram_r_3_6_port, d => 
                           n528, outb => n1297);
   U1801 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_7_6_port, b
                           => n529, outb => n1296);
   U1802 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_1_6_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_0_block_ram_r_0_6_port, d => 
                           n531, outb => n1295);
   U1803 : aoi22 port map( a => n532, b => n1209, c => n534, d => n1223, outb 
                           => n1293);
   U1804 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_2_6_port, 
                           outb => n1223);
   U1805 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_4_6_port, 
                           outb => n1209);
   U1806 : nand2 port map( a => n536, b => n1195, outb => n1292);
   U1807 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_6_6_port, 
                           outb => n1195);
   U1808 : nand4 port map( a => n538, b => n1298, c => n1299, d => n1300, outb 
                           => n1289);
   U1809 : nor3 port map( a => n1301, b => n1302, c => n1303, outb => n1300);
   U1810 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_13_6_port,
                           b => n527, c => 
                           load_n_store_RGB_Array_0_block_ram_r_11_6_port, d =>
                           n528, outb => n1303);
   U1811 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_15_6_port, 
                           b => n529, outb => n1302);
   U1812 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_9_6_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_0_block_ram_r_8_6_port, d => 
                           n531, outb => n1301);
   U1813 : aoi22 port map( a => n532, b => n1147, c => n534, d => n1162, outb 
                           => n1299);
   U1814 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_10_6_port,
                           outb => n1162);
   U1815 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_12_6_port,
                           outb => n1147);
   U1816 : nand2 port map( a => n536, b => n1105, outb => n1298);
   U1817 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_14_6_port,
                           outb => n1105);
   U1818 : nand3 port map( a => n1304, b => n1305, c => n1306, outb => 
                           load_n_store_RGB_Array_0_n128);
   U1819 : nand2 port map( a => load_n_store_lazy_in_0_5_port, b => 
                           load_n_store_we_i, outb => n1306);
   U1820 : nand4 port map( a => n520, b => n1307, c => n1308, d => n1309, outb 
                           => n1305);
   U1821 : nor3 port map( a => n1310, b => n1311, c => n1312, outb => n1309);
   U1822 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_5_5_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_0_block_ram_r_3_5_port, d => 
                           n528, outb => n1312);
   U1823 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_7_5_port, b
                           => n529, outb => n1311);
   U1824 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_1_5_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_0_block_ram_r_0_5_port, d => 
                           n531, outb => n1310);
   U1825 : aoi22 port map( a => n532, b => n1210, c => n534, d => n1224, outb 
                           => n1308);
   U1826 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_2_5_port, 
                           outb => n1224);
   U1827 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_4_5_port, 
                           outb => n1210);
   U1828 : nand2 port map( a => n536, b => n1196, outb => n1307);
   U1829 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_6_5_port, 
                           outb => n1196);
   U1830 : nand4 port map( a => n538, b => n1313, c => n1314, d => n1315, outb 
                           => n1304);
   U1831 : nor3 port map( a => n1316, b => n1317, c => n1318, outb => n1315);
   U1832 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_13_5_port,
                           b => n527, c => 
                           load_n_store_RGB_Array_0_block_ram_r_11_5_port, d =>
                           n528, outb => n1318);
   U1833 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_15_5_port, 
                           b => n529, outb => n1317);
   U1834 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_9_5_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_0_block_ram_r_8_5_port, d => 
                           n531, outb => n1316);
   U1835 : aoi22 port map( a => n532, b => n1148, c => n534, d => n1163, outb 
                           => n1314);
   U1836 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_10_5_port,
                           outb => n1163);
   U1837 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_12_5_port,
                           outb => n1148);
   U1838 : nand2 port map( a => n536, b => n1107, outb => n1313);
   U1839 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_14_5_port,
                           outb => n1107);
   U1840 : nand3 port map( a => n1319, b => n1320, c => n1321, outb => 
                           load_n_store_RGB_Array_0_n105);
   U1841 : nand2 port map( a => load_n_store_lazy_in_0_4_port, b => 
                           load_n_store_we_i, outb => n1321);
   U1842 : nand4 port map( a => n520, b => n1322, c => n1323, d => n1324, outb 
                           => n1320);
   U1843 : nor3 port map( a => n1325, b => n1326, c => n1327, outb => n1324);
   U1844 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_5_4_port, 
                           b => n527, c => 
                           load_n_store_RGB_Array_0_block_ram_r_3_4_port, d => 
                           n528, outb => n1327);
   U1845 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_7_4_port, b
                           => n529, outb => n1326);
   U1846 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_1_4_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_0_block_ram_r_0_4_port, d => 
                           n531, outb => n1325);
   U1847 : aoi22 port map( a => n532, b => n1211, c => n534, d => n1225, outb 
                           => n1323);
   U1848 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_2_4_port, 
                           outb => n1225);
   U1849 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_4_4_port, 
                           outb => n1211);
   U1850 : nand2 port map( a => n536, b => n1197, outb => n1322);
   U1851 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_6_4_port, 
                           outb => n1197);
   U1852 : nor2 port map( a => addr_i_3_port, b => load_n_store_we_i, outb => 
                           n520);
   U1853 : nand4 port map( a => n538, b => n1328, c => n1329, d => n1330, outb 
                           => n1319);
   U1854 : nor3 port map( a => n1331, b => n1332, c => n1333, outb => n1330);
   U1855 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_13_4_port,
                           b => n527, c => 
                           load_n_store_RGB_Array_0_block_ram_r_11_4_port, d =>
                           n528, outb => n1333);
   U1856 : inv port map( inb => n1160, outb => n528);
   U1857 : nor3 port map( a => n20, b => addr_i_2_port, c => n24, outb => n1160
                           );
   U1858 : inv port map( inb => n1145, outb => n527);
   U1859 : nor3 port map( a => n24, b => addr_i_1_port, c => n52, outb => n1145
                           );
   U1860 : nor2 port map( a => load_n_store_RGB_Array_0_block_ram_r_15_4_port, 
                           b => n529, outb => n1332);
   U1861 : inv port map( inb => n1101, outb => n529);
   U1862 : nor3 port map( a => n24, b => n20, c => n52, outb => n1101);
   U1863 : oai22 port map( a => load_n_store_RGB_Array_0_block_ram_r_9_4_port, 
                           b => n530, c => 
                           load_n_store_RGB_Array_0_block_ram_r_8_4_port, d => 
                           n531, outb => n1331);
   U1864 : inv port map( inb => n1184, outb => n531);
   U1865 : nor3 port map( a => addr_i_1_port, b => addr_i_2_port, c => 
                           addr_i_0_port, outb => n1184);
   U1866 : inv port map( inb => n1175, outb => n530);
   U1867 : nor3 port map( a => addr_i_1_port, b => addr_i_2_port, c => n24, 
                           outb => n1175);
   U1868 : inv port map( inb => addr_i_0_port, outb => n24);
   U1869 : aoi22 port map( a => n532, b => n1149, c => n534, d => n1164, outb 
                           => n1329);
   U1870 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_10_4_port,
                           outb => n1164);
   U1871 : nor3 port map( a => addr_i_0_port, b => addr_i_2_port, c => n20, 
                           outb => n534);
   U1872 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_12_4_port,
                           outb => n1149);
   U1873 : nor3 port map( a => addr_i_0_port, b => addr_i_1_port, c => n52, 
                           outb => n532);
   U1874 : nand2 port map( a => n536, b => n1130, outb => n1328);
   U1875 : inv port map( inb => load_n_store_RGB_Array_0_block_ram_r_14_4_port,
                           outb => n1130);
   U1876 : nor3 port map( a => n20, b => addr_i_0_port, c => n52, outb => n536)
                           ;
   U1877 : inv port map( inb => addr_i_2_port, outb => n52);
   U1878 : inv port map( inb => addr_i_1_port, outb => n20);
   U1879 : nor2 port map( a => n46, b => load_n_store_we_i, outb => n538);
   U1880 : inv port map( inb => addr_i_3_port, outb => n46);
   U1881 : oai12 port map( b => n1334, c => n1335, a => n1336, outb => 
                           display_out_n912);
   U1882 : nand2 port map( a => n1337, b => n1335, outb => n1336);
   U1883 : nand4 port map( a => n1338, b => n1339, c => n1340, d => n1341, outb
                           => n1337);
   U1884 : aoi22 port map( a => n1342, b => n1343, c => n1344, d => n1345, outb
                           => n1341);
   U1885 : nand2 port map( a => n1346, b => reg_hub_f, outb => n1340);
   U1886 : oai22 port map( a => n1347, b => n1348, c => n1349, d => n1335, outb
                           => display_out_n911);
   U1887 : nor2 port map( a => n1350, b => n1351, outb => n1348);
   U1888 : nor3 port map( a => n1352, b => reg_hub_f, c => n501, outb => n1351)
                           ;
   U1889 : oai22 port map( a => n1353, b => n1354, c => n1355, d => n402, outb 
                           => display_out_n910);
   U1890 : inv port map( inb => display_out_clk_timer_31_port, outb => n1353);
   U1891 : oai22 port map( a => n1356, b => n1357, c => n402, d => n1358, outb 
                           => display_out_n909);
   U1892 : xor2 port map( a => n1359, b => n1360, outb => n402);
   U1893 : aoi22 port map( a => n1361, b => n1362, c => n1363, d => n1364, outb
                           => n1360);
   U1894 : inv port map( inb => n1365, outb => n1362);
   U1895 : nor2 port map( a => n1364, b => n1363, outb => n1365);
   U1896 : xor2 port map( a => n1366, b => n1361, outb => n1359);
   U1897 : oai12 port map( b => n1356, c => n1367, a => n1368, outb => n1366);
   U1898 : aoi22 port map( a => display_out_clk_timer_31_port, b => n1369, c =>
                           display_out_h_row_31_port, d => n1370, outb => n1368
                           );
   U1899 : inv port map( inb => display_out_h_col_31_port, outb => n1356);
   U1900 : oai22 port map( a => n1371, b => n1372, c => n1373, d => n1354, outb
                           => display_out_n908);
   U1901 : aoi12 port map( b => n422, c => n1374, a => n1375, outb => n1372);
   U1902 : inv port map( inb => n1376, outb => n1375);
   U1903 : oai22 port map( a => n1377, b => n1354, c => n1355, d => n400, outb 
                           => display_out_n907);
   U1904 : oai22 port map( a => n1378, b => n1354, c => n1355, d => n398, outb 
                           => display_out_n906);
   U1905 : oai22 port map( a => n1379, b => n1354, c => n1355, d => n396, outb 
                           => display_out_n905);
   U1906 : oai22 port map( a => n1380, b => n1354, c => n1355, d => n394, outb 
                           => display_out_n904);
   U1907 : oai22 port map( a => n1381, b => n1354, c => n1355, d => n392, outb 
                           => display_out_n903);
   U1908 : oai22 port map( a => n1382, b => n1354, c => n1355, d => n390, outb 
                           => display_out_n902);
   U1909 : oai22 port map( a => n1383, b => n1354, c => n1355, d => n388, outb 
                           => display_out_n901);
   U1910 : oai22 port map( a => n1384, b => n1354, c => n1355, d => n386, outb 
                           => display_out_n900);
   U1911 : oai22 port map( a => n1385, b => n1354, c => n1355, d => n384, outb 
                           => display_out_n899);
   U1912 : oai22 port map( a => n1386, b => n1354, c => n1355, d => n382, outb 
                           => display_out_n898);
   U1913 : oai22 port map( a => n1387, b => n1354, c => n1355, d => n380, outb 
                           => display_out_n897);
   U1914 : oai22 port map( a => n1388, b => n1354, c => n1355, d => n378, outb 
                           => display_out_n896);
   U1915 : oai22 port map( a => n1389, b => n1354, c => n1355, d => n376, outb 
                           => display_out_n895);
   U1916 : oai22 port map( a => n1390, b => n1354, c => n1355, d => n374, outb 
                           => display_out_n894);
   U1917 : oai22 port map( a => n1391, b => n1354, c => n1355, d => n372, outb 
                           => display_out_n893);
   U1918 : oai22 port map( a => n1392, b => n1354, c => n1355, d => n370, outb 
                           => display_out_n892);
   U1919 : inv port map( inb => display_out_clk_timer_15_port, outb => n1392);
   U1920 : oai22 port map( a => n1393, b => n1354, c => n1355, d => n368, outb 
                           => display_out_n891);
   U1921 : inv port map( inb => display_out_clk_timer_14_port, outb => n1393);
   U1922 : oai22 port map( a => n1394, b => n1354, c => n1355, d => n366, outb 
                           => display_out_n890);
   U1923 : inv port map( inb => display_out_clk_timer_13_port, outb => n1394);
   U1924 : oai22 port map( a => n1395, b => n1354, c => n1355, d => n364, outb 
                           => display_out_n889);
   U1925 : inv port map( inb => display_out_clk_timer_12_port, outb => n1395);
   U1926 : oai22 port map( a => n1396, b => n1354, c => n1355, d => n362, outb 
                           => display_out_n888);
   U1927 : inv port map( inb => display_out_clk_timer_11_port, outb => n1396);
   U1928 : oai22 port map( a => n1397, b => n1354, c => n1355, d => n359, outb 
                           => display_out_n887);
   U1929 : inv port map( inb => display_out_clk_timer_10_port, outb => n1397);
   U1930 : oai22 port map( a => n1398, b => n1354, c => n1355, d => n404, outb 
                           => display_out_n886);
   U1931 : oai22 port map( a => n1399, b => n1354, c => n1355, d => n406, outb 
                           => display_out_n885);
   U1932 : oai22 port map( a => n1400, b => n1354, c => n1355, d => n408, outb 
                           => display_out_n884);
   U1933 : oai22 port map( a => n1401, b => n1354, c => n1355, d => n410, outb 
                           => display_out_n883);
   U1934 : oai22 port map( a => n1402, b => n1354, c => n1355, d => n412, outb 
                           => display_out_n882);
   U1935 : oai12 port map( b => n1355, c => n414, a => n1403, outb => 
                           display_out_n881);
   U1936 : aoi22 port map( a => n1404, b => n1354, c => n1371, d => 
                           display_out_clk_timer_4_port, outb => n1403);
   U1937 : nand2 port map( a => n1405, b => n1376, outb => display_out_n880);
   U1938 : nor2 port map( a => n1346, b => n1406, outb => n1376);
   U1939 : aoi22 port map( a => n417, b => n1374, c => n1371, d => 
                           display_out_clk_timer_3_port, outb => n1405);
   U1940 : inv port map( inb => n1407, outb => n417);
   U1941 : oai12 port map( b => n1355, c => n420, a => n1408, outb => 
                           display_out_n879);
   U1942 : aoi22 port map( a => n1404, b => n1354, c => n1371, d => 
                           display_out_clk_timer_2_port, outb => n1408);
   U1943 : inv port map( inb => n1354, outb => n1371);
   U1944 : oai22 port map( a => n1409, b => n1354, c => n1355, d => n424, outb 
                           => display_out_n878);
   U1945 : inv port map( inb => n1410, outb => n1355);
   U1946 : nand4 port map( a => n1411, b => n1412, c => n1413, d => n1414, outb
                           => n1354);
   U1947 : inv port map( inb => display_out_clk_timer_1_port, outb => n1409);
   U1948 : nand4 port map( a => n1415, b => n1416, c => n1417, d => n1339, outb
                           => display_out_n877);
   U1949 : nand2 port map( a => n1347, b => display_out_hub_out_sm_1_port, outb
                           => n1417);
   U1950 : inv port map( inb => n1335, outb => n1347);
   U1951 : nand4 port map( a => n1418, b => n1419, c => n1420, d => n1421, outb
                           => n1335);
   U1952 : nand2 port map( a => n1346, b => mem_hub_f, outb => n1420);
   U1953 : nand2 port map( a => n1342, b => n1422, outb => n1416);
   U1954 : oai22 port map( a => n1423, b => n1357, c => n1424, d => n1358, outb
                           => display_out_n876);
   U1955 : oai22 port map( a => n1425, b => n1357, c => n400, d => n1358, outb 
                           => display_out_n875);
   U1956 : xor2 port map( a => n1363, b => n1426, outb => n400);
   U1957 : xor2 port map( a => n1361, b => n1364, outb => n1426);
   U1958 : inv port map( inb => n1427, outb => n1364);
   U1959 : oai12 port map( b => n1367, c => n1425, a => n1428, outb => n1427);
   U1960 : aoi22 port map( a => display_out_clk_timer_30_port, b => n1369, c =>
                           display_out_h_row_30_port, d => n1370, outb => n1428
                           );
   U1961 : aoi22 port map( a => n1429, b => n1430, c => n1369, d => n1431, outb
                           => n1363);
   U1962 : inv port map( inb => n1432, outb => n1431);
   U1963 : nor2 port map( a => n1430, b => n1429, outb => n1432);
   U1964 : oai22 port map( a => n1433, b => n1357, c => n398, d => n1358, outb 
                           => display_out_n874);
   U1965 : xor2 port map( a => n1434, b => n1430, outb => n398);
   U1966 : aoi22 port map( a => n1435, b => n1436, c => n1437, d => n1361, outb
                           => n1430);
   U1967 : inv port map( inb => n1438, outb => n1437);
   U1968 : nor2 port map( a => n1436, b => n1435, outb => n1438);
   U1969 : xor2 port map( a => n1429, b => n1361, outb => n1434);
   U1970 : oai12 port map( b => n1367, c => n1433, a => n1439, outb => n1429);
   U1971 : aoi22 port map( a => display_out_clk_timer_29_port, b => n1369, c =>
                           display_out_h_row_29_port, d => n1370, outb => n1439
                           );
   U1972 : oai22 port map( a => n1440, b => n1357, c => n396, d => n1358, outb 
                           => display_out_n873);
   U1973 : xor2 port map( a => n1436, b => n1441, outb => n396);
   U1974 : xor2 port map( a => n1361, b => n1435, outb => n1441);
   U1975 : inv port map( inb => n1442, outb => n1435);
   U1976 : oai12 port map( b => n1367, c => n1440, a => n1443, outb => n1442);
   U1977 : aoi22 port map( a => display_out_clk_timer_28_port, b => n1369, c =>
                           display_out_h_row_28_port, d => n1370, outb => n1443
                           );
   U1978 : aoi22 port map( a => n1444, b => n1445, c => n1369, d => n1446, outb
                           => n1436);
   U1979 : inv port map( inb => n1447, outb => n1446);
   U1980 : nor2 port map( a => n1445, b => n1444, outb => n1447);
   U1981 : oai22 port map( a => n1448, b => n1357, c => n394, d => n1358, outb 
                           => display_out_n872);
   U1982 : xor2 port map( a => n1449, b => n1445, outb => n394);
   U1983 : aoi22 port map( a => n1450, b => n1451, c => n1452, d => n1361, outb
                           => n1445);
   U1984 : inv port map( inb => n1453, outb => n1452);
   U1985 : nor2 port map( a => n1451, b => n1450, outb => n1453);
   U1986 : xor2 port map( a => n1444, b => n1361, outb => n1449);
   U1987 : oai12 port map( b => n1367, c => n1448, a => n1454, outb => n1444);
   U1988 : aoi22 port map( a => display_out_clk_timer_27_port, b => n1369, c =>
                           display_out_h_row_27_port, d => n1370, outb => n1454
                           );
   U1989 : oai22 port map( a => n1455, b => n1357, c => n392, d => n1358, outb 
                           => display_out_n871);
   U1990 : xor2 port map( a => n1451, b => n1456, outb => n392);
   U1991 : xor2 port map( a => n1361, b => n1450, outb => n1456);
   U1992 : inv port map( inb => n1457, outb => n1450);
   U1993 : oai12 port map( b => n1367, c => n1455, a => n1458, outb => n1457);
   U1994 : aoi22 port map( a => display_out_clk_timer_26_port, b => n1369, c =>
                           display_out_h_row_26_port, d => n1370, outb => n1458
                           );
   U1995 : aoi22 port map( a => n1459, b => n1460, c => n1369, d => n1461, outb
                           => n1451);
   U1996 : inv port map( inb => n1462, outb => n1461);
   U1997 : nor2 port map( a => n1460, b => n1459, outb => n1462);
   U1998 : oai22 port map( a => n1463, b => n1357, c => n390, d => n1358, outb 
                           => display_out_n870);
   U1999 : xor2 port map( a => n1464, b => n1460, outb => n390);
   U2000 : aoi22 port map( a => n1465, b => n1466, c => n1467, d => n1361, outb
                           => n1460);
   U2001 : nand2 port map( a => n1468, b => n1469, outb => n1467);
   U2002 : xor2 port map( a => n1459, b => n1361, outb => n1464);
   U2003 : oai12 port map( b => n1367, c => n1463, a => n1470, outb => n1459);
   U2004 : aoi22 port map( a => display_out_clk_timer_25_port, b => n1369, c =>
                           display_out_h_row_25_port, d => n1370, outb => n1470
                           );
   U2005 : oai22 port map( a => n1471, b => n1357, c => n388, d => n1358, outb 
                           => display_out_n869);
   U2006 : xor2 port map( a => n1472, b => n1469, outb => n388);
   U2007 : inv port map( inb => n1465, outb => n1469);
   U2008 : oai22 port map( a => n1473, b => n1474, c => n1475, d => n1369, outb
                           => n1465);
   U2009 : inv port map( inb => n1476, outb => n1475);
   U2010 : nand2 port map( a => n1474, b => n1473, outb => n1476);
   U2011 : xor2 port map( a => n1466, b => n1369, outb => n1472);
   U2012 : inv port map( inb => n1468, outb => n1466);
   U2013 : oai12 port map( b => n1367, c => n1471, a => n1477, outb => n1468);
   U2014 : aoi22 port map( a => display_out_clk_timer_24_port, b => n1369, c =>
                           display_out_h_row_24_port, d => n1370, outb => n1477
                           );
   U2015 : oai22 port map( a => n1478, b => n1357, c => n386, d => n1358, outb 
                           => display_out_n868);
   U2016 : xor2 port map( a => n1479, b => n1473, outb => n386);
   U2017 : aoi22 port map( a => n1480, b => n1481, c => n1482, d => n1361, outb
                           => n1473);
   U2018 : nand2 port map( a => n1483, b => n1484, outb => n1482);
   U2019 : inv port map( inb => n1483, outb => n1481);
   U2020 : xor2 port map( a => n1474, b => n1361, outb => n1479);
   U2021 : oai12 port map( b => n1367, c => n1478, a => n1485, outb => n1474);
   U2022 : aoi22 port map( a => display_out_clk_timer_23_port, b => n1369, c =>
                           display_out_h_row_23_port, d => n1370, outb => n1485
                           );
   U2023 : oai22 port map( a => n1486, b => n1357, c => n384, d => n1358, outb 
                           => display_out_n867);
   U2024 : xor2 port map( a => n1487, b => n1484, outb => n384);
   U2025 : inv port map( inb => n1480, outb => n1484);
   U2026 : oai22 port map( a => n1488, b => n1489, c => n1490, d => n1369, outb
                           => n1480);
   U2027 : inv port map( inb => n1491, outb => n1490);
   U2028 : nand2 port map( a => n1489, b => n1488, outb => n1491);
   U2029 : xor2 port map( a => n1483, b => n1361, outb => n1487);
   U2030 : oai12 port map( b => n1367, c => n1486, a => n1492, outb => n1483);
   U2031 : aoi22 port map( a => display_out_clk_timer_22_port, b => n1369, c =>
                           display_out_h_row_22_port, d => n1370, outb => n1492
                           );
   U2032 : oai22 port map( a => n1493, b => n1357, c => n382, d => n1358, outb 
                           => display_out_n866);
   U2033 : xor2 port map( a => n1494, b => n1488, outb => n382);
   U2034 : aoi22 port map( a => n1495, b => n1496, c => n1497, d => n1361, outb
                           => n1488);
   U2035 : nand2 port map( a => n1498, b => n1499, outb => n1497);
   U2036 : inv port map( inb => n1498, outb => n1496);
   U2037 : xor2 port map( a => n1489, b => n1361, outb => n1494);
   U2038 : oai12 port map( b => n1367, c => n1493, a => n1500, outb => n1489);
   U2039 : aoi22 port map( a => display_out_clk_timer_21_port, b => n1369, c =>
                           display_out_h_row_21_port, d => n1370, outb => n1500
                           );
   U2040 : oai22 port map( a => n1501, b => n1357, c => n380, d => n1358, outb 
                           => display_out_n865);
   U2041 : xor2 port map( a => n1502, b => n1499, outb => n380);
   U2042 : inv port map( inb => n1495, outb => n1499);
   U2043 : oai22 port map( a => n1503, b => n1504, c => n1505, d => n1369, outb
                           => n1495);
   U2044 : inv port map( inb => n1506, outb => n1505);
   U2045 : nand2 port map( a => n1504, b => n1503, outb => n1506);
   U2046 : xor2 port map( a => n1498, b => n1361, outb => n1502);
   U2047 : oai12 port map( b => n1367, c => n1501, a => n1507, outb => n1498);
   U2048 : aoi22 port map( a => display_out_clk_timer_20_port, b => n1369, c =>
                           display_out_h_row_20_port, d => n1370, outb => n1507
                           );
   U2049 : oai22 port map( a => n1508, b => n1357, c => n378, d => n1358, outb 
                           => display_out_n864);
   U2050 : xor2 port map( a => n1509, b => n1503, outb => n378);
   U2051 : aoi22 port map( a => n1510, b => n1511, c => n1512, d => n1361, outb
                           => n1503);
   U2052 : nand2 port map( a => n1513, b => n1514, outb => n1512);
   U2053 : inv port map( inb => n1513, outb => n1511);
   U2054 : xor2 port map( a => n1504, b => n1361, outb => n1509);
   U2055 : oai12 port map( b => n1367, c => n1508, a => n1515, outb => n1504);
   U2056 : aoi22 port map( a => display_out_clk_timer_19_port, b => n1369, c =>
                           display_out_h_row_19_port, d => n1370, outb => n1515
                           );
   U2057 : oai22 port map( a => n1516, b => n1357, c => n376, d => n1358, outb 
                           => display_out_n863);
   U2058 : xor2 port map( a => n1517, b => n1514, outb => n376);
   U2059 : inv port map( inb => n1510, outb => n1514);
   U2060 : oai22 port map( a => n1518, b => n1519, c => n1520, d => n1369, outb
                           => n1510);
   U2061 : inv port map( inb => n1521, outb => n1520);
   U2062 : nand2 port map( a => n1519, b => n1518, outb => n1521);
   U2063 : xor2 port map( a => n1513, b => n1361, outb => n1517);
   U2064 : oai12 port map( b => n1367, c => n1516, a => n1522, outb => n1513);
   U2065 : aoi22 port map( a => display_out_clk_timer_18_port, b => n1369, c =>
                           display_out_h_row_18_port, d => n1370, outb => n1522
                           );
   U2066 : oai22 port map( a => n1523, b => n1357, c => n374, d => n1358, outb 
                           => display_out_n862);
   U2067 : xor2 port map( a => n1524, b => n1518, outb => n374);
   U2068 : aoi22 port map( a => n1525, b => n1526, c => n1527, d => n1361, outb
                           => n1518);
   U2069 : nand2 port map( a => n1528, b => n1529, outb => n1527);
   U2070 : inv port map( inb => n1528, outb => n1526);
   U2071 : xor2 port map( a => n1519, b => n1361, outb => n1524);
   U2072 : oai12 port map( b => n1367, c => n1523, a => n1530, outb => n1519);
   U2073 : aoi22 port map( a => display_out_clk_timer_17_port, b => n1369, c =>
                           display_out_h_row_17_port, d => n1370, outb => n1530
                           );
   U2074 : oai22 port map( a => n1531, b => n1357, c => n372, d => n1358, outb 
                           => display_out_n861);
   U2075 : xor2 port map( a => n1532, b => n1529, outb => n372);
   U2076 : inv port map( inb => n1525, outb => n1529);
   U2077 : oai22 port map( a => n1533, b => n1534, c => n1535, d => n1369, outb
                           => n1525);
   U2078 : inv port map( inb => n1536, outb => n1535);
   U2079 : nand2 port map( a => n1534, b => n1533, outb => n1536);
   U2080 : xor2 port map( a => n1528, b => n1361, outb => n1532);
   U2081 : oai12 port map( b => n1367, c => n1531, a => n1537, outb => n1528);
   U2082 : aoi22 port map( a => display_out_clk_timer_16_port, b => n1369, c =>
                           display_out_h_row_16_port, d => n1370, outb => n1537
                           );
   U2083 : oai22 port map( a => n1538, b => n1357, c => n370, d => n1358, outb 
                           => display_out_n860);
   U2084 : xor2 port map( a => n1539, b => n1533, outb => n370);
   U2085 : aoi22 port map( a => n1540, b => n1541, c => n1542, d => n1361, outb
                           => n1533);
   U2086 : nand2 port map( a => n1543, b => n1544, outb => n1542);
   U2087 : inv port map( inb => n1543, outb => n1541);
   U2088 : xor2 port map( a => n1534, b => n1361, outb => n1539);
   U2089 : oai12 port map( b => n1367, c => n1538, a => n1545, outb => n1534);
   U2090 : aoi22 port map( a => display_out_clk_timer_15_port, b => n1369, c =>
                           display_out_h_row_15_port, d => n1370, outb => n1545
                           );
   U2091 : oai22 port map( a => n1546, b => n1357, c => n368, d => n1358, outb 
                           => display_out_n859);
   U2092 : xor2 port map( a => n1547, b => n1544, outb => n368);
   U2093 : inv port map( inb => n1540, outb => n1544);
   U2094 : oai22 port map( a => n1548, b => n1549, c => n1550, d => n1369, outb
                           => n1540);
   U2095 : inv port map( inb => n1551, outb => n1550);
   U2096 : nand2 port map( a => n1549, b => n1548, outb => n1551);
   U2097 : xor2 port map( a => n1543, b => n1361, outb => n1547);
   U2098 : oai12 port map( b => n1367, c => n1546, a => n1552, outb => n1543);
   U2099 : aoi22 port map( a => display_out_clk_timer_14_port, b => n1369, c =>
                           display_out_h_row_14_port, d => n1370, outb => n1552
                           );
   U2100 : oai22 port map( a => n1553, b => n1357, c => n366, d => n1358, outb 
                           => display_out_n858);
   U2101 : xor2 port map( a => n1554, b => n1548, outb => n366);
   U2102 : aoi22 port map( a => n1555, b => n1556, c => n1557, d => n1361, outb
                           => n1548);
   U2103 : nand2 port map( a => n1558, b => n1559, outb => n1557);
   U2104 : inv port map( inb => n1558, outb => n1556);
   U2105 : xor2 port map( a => n1549, b => n1361, outb => n1554);
   U2106 : oai12 port map( b => n1367, c => n1553, a => n1560, outb => n1549);
   U2107 : aoi22 port map( a => display_out_clk_timer_13_port, b => n1369, c =>
                           display_out_h_row_13_port, d => n1370, outb => n1560
                           );
   U2108 : oai22 port map( a => n1561, b => n1357, c => n364, d => n1358, outb 
                           => display_out_n857);
   U2109 : xor2 port map( a => n1562, b => n1559, outb => n364);
   U2110 : inv port map( inb => n1555, outb => n1559);
   U2111 : oai22 port map( a => n1563, b => n1564, c => n1565, d => n1369, outb
                           => n1555);
   U2112 : inv port map( inb => n1566, outb => n1565);
   U2113 : nand2 port map( a => n1564, b => n1563, outb => n1566);
   U2114 : xor2 port map( a => n1558, b => n1361, outb => n1562);
   U2115 : oai12 port map( b => n1367, c => n1561, a => n1567, outb => n1558);
   U2116 : aoi22 port map( a => display_out_clk_timer_12_port, b => n1369, c =>
                           display_out_h_row_12_port, d => n1370, outb => n1567
                           );
   U2117 : oai22 port map( a => n1568, b => n1357, c => n362, d => n1358, outb 
                           => display_out_n856);
   U2118 : xor2 port map( a => n1569, b => n1564, outb => n362);
   U2119 : oai12 port map( b => n1367, c => n1568, a => n1570, outb => n1564);
   U2120 : aoi22 port map( a => display_out_clk_timer_11_port, b => n1369, c =>
                           display_out_h_row_11_port, d => n1370, outb => n1570
                           );
   U2121 : xor2 port map( a => n1563, b => n1361, outb => n1569);
   U2122 : oai22 port map( a => n1571, b => n1572, c => n1361, d => n1573, outb
                           => n1563);
   U2123 : inv port map( inb => n1574, outb => n1573);
   U2124 : nand2 port map( a => n1572, b => n1571, outb => n1574);
   U2125 : oai22 port map( a => n1575, b => n1357, c => n359, d => n1358, outb 
                           => display_out_n855);
   U2126 : xor2 port map( a => n1576, b => n1571, outb => n359);
   U2127 : inv port map( inb => n1577, outb => n1571);
   U2128 : oai12 port map( b => n1367, c => n1575, a => n1578, outb => n1577);
   U2129 : aoi22 port map( a => display_out_clk_timer_10_port, b => n1369, c =>
                           display_out_h_row_10_port, d => n1370, outb => n1578
                           );
   U2130 : xor2 port map( a => n1361, b => n1572, outb => n1576);
   U2131 : oai22 port map( a => n1579, b => n1580, c => n1581, d => n1369, outb
                           => n1572);
   U2132 : inv port map( inb => n1582, outb => n1581);
   U2133 : nand2 port map( a => n1579, b => n1580, outb => n1582);
   U2134 : oai22 port map( a => n1583, b => n1357, c => n404, d => n1358, outb 
                           => display_out_n854);
   U2135 : xor2 port map( a => n1584, b => n1579, outb => n404);
   U2136 : oai12 port map( b => n1367, c => n1583, a => n1585, outb => n1579);
   U2137 : aoi22 port map( a => display_out_clk_timer_9_port, b => n1369, c => 
                           display_out_h_row_9_port, d => n1370, outb => n1585)
                           ;
   U2138 : xor2 port map( a => n1580, b => n1361, outb => n1584);
   U2139 : oai22 port map( a => n1586, b => n1587, c => n1361, d => n1588, outb
                           => n1580);
   U2140 : inv port map( inb => n1589, outb => n1588);
   U2141 : nand2 port map( a => n1587, b => n1586, outb => n1589);
   U2142 : oai22 port map( a => n1590, b => n1357, c => n406, d => n1358, outb 
                           => display_out_n853);
   U2143 : xor2 port map( a => n1591, b => n1586, outb => n406);
   U2144 : inv port map( inb => n1592, outb => n1586);
   U2145 : oai12 port map( b => n1367, c => n1590, a => n1593, outb => n1592);
   U2146 : aoi22 port map( a => display_out_clk_timer_8_port, b => n1369, c => 
                           display_out_h_row_8_port, d => n1370, outb => n1593)
                           ;
   U2147 : xor2 port map( a => n1361, b => n1587, outb => n1591);
   U2148 : oai22 port map( a => n1594, b => n1595, c => n1596, d => n1369, outb
                           => n1587);
   U2149 : nor2 port map( a => n1597, b => n1598, outb => n1596);
   U2150 : inv port map( inb => n1594, outb => n1597);
   U2151 : inv port map( inb => n1598, outb => n1595);
   U2152 : oai22 port map( a => n1599, b => n1357, c => n408, d => n1358, outb 
                           => display_out_n852);
   U2153 : xor2 port map( a => n1600, b => n1594, outb => n408);
   U2154 : oai12 port map( b => n1367, c => n1599, a => n1601, outb => n1594);
   U2155 : aoi22 port map( a => display_out_clk_timer_7_port, b => n1369, c => 
                           display_out_h_row_7_port, d => n1370, outb => n1601)
                           ;
   U2156 : xor2 port map( a => n1598, b => n1369, outb => n1600);
   U2157 : aoi22 port map( a => n1602, b => n1603, c => n1369, d => n1604, outb
                           => n1598);
   U2158 : inv port map( inb => n1605, outb => n1604);
   U2159 : nor2 port map( a => n1603, b => n1602, outb => n1605);
   U2160 : oai22 port map( a => n1606, b => n1357, c => n410, d => n1358, outb 
                           => display_out_n851);
   U2161 : xor2 port map( a => n1607, b => n1603, outb => n410);
   U2162 : oai12 port map( b => n1367, c => n1606, a => n1608, outb => n1603);
   U2163 : aoi22 port map( a => display_out_clk_timer_6_port, b => n1369, c => 
                           display_out_h_row_6_port, d => n1370, outb => n1608)
                           ;
   U2164 : xor2 port map( a => n1602, b => n1361, outb => n1607);
   U2165 : oai22 port map( a => n1609, b => n1610, c => n1361, d => n1611, outb
                           => n1602);
   U2166 : inv port map( inb => n1612, outb => n1611);
   U2167 : nand2 port map( a => n1610, b => n1609, outb => n1612);
   U2168 : oai22 port map( a => n1613, b => n1357, c => n412, d => n1358, outb 
                           => display_out_n850);
   U2169 : xor2 port map( a => n1614, b => n1609, outb => n412);
   U2170 : inv port map( inb => n1615, outb => n1609);
   U2171 : oai12 port map( b => n1367, c => n1613, a => n1616, outb => n1615);
   U2172 : aoi22 port map( a => display_out_clk_timer_5_port, b => n1369, c => 
                           display_out_h_row_5_port, d => n1370, outb => n1616)
                           ;
   U2173 : xor2 port map( a => n1361, b => n1610, outb => n1614);
   U2174 : oai22 port map( a => n1617, b => n1618, c => n1619, d => n1369, outb
                           => n1610);
   U2175 : inv port map( inb => n1620, outb => n1619);
   U2176 : nand2 port map( a => n1617, b => n1618, outb => n1620);
   U2177 : oai22 port map( a => n1621, b => n1357, c => n414, d => n1358, outb 
                           => display_out_n849);
   U2178 : xor2 port map( a => n1622, b => n1617, outb => n414);
   U2179 : oai12 port map( b => n1367, c => n1621, a => n1623, outb => n1617);
   U2180 : aoi22 port map( a => display_out_clk_timer_4_port, b => n1369, c => 
                           display_out_h_row_4_port, d => n1370, outb => n1623)
                           ;
   U2181 : xor2 port map( a => n1618, b => n1361, outb => n1622);
   U2182 : oai22 port map( a => n1624, b => n1625, c => n1361, d => n1626, outb
                           => n1618);
   U2183 : nor2 port map( a => n1627, b => n1628, outb => n1626);
   U2184 : inv port map( inb => n1628, outb => n1624);
   U2185 : oai22 port map( a => n1629, b => n1357, c => n1407, d => n1358, outb
                           => display_out_n848);
   U2186 : xor2 port map( a => n1630, b => n1627, outb => n1407);
   U2187 : inv port map( inb => n1625, outb => n1627);
   U2188 : oai22 port map( a => n1631, b => n1632, c => n1633, d => n1369, outb
                           => n1625);
   U2189 : inv port map( inb => n1634, outb => n1633);
   U2190 : nand2 port map( a => n1632, b => n1631, outb => n1634);
   U2191 : xor2 port map( a => n1628, b => n1361, outb => n1630);
   U2192 : oai12 port map( b => n1367, c => n1629, a => n1635, outb => n1628);
   U2193 : aoi22 port map( a => display_out_clk_timer_3_port, b => n1369, c => 
                           display_out_h_row_3_port, d => n1370, outb => n1635)
                           ;
   U2194 : oai22 port map( a => n1636, b => n1357, c => n420, d => n1358, outb 
                           => display_out_n847);
   U2195 : xor2 port map( a => n1637, b => n1631, outb => n420);
   U2196 : aoi22 port map( a => n1638, b => n422, c => n1639, d => n1361, outb 
                           => n1631);
   U2197 : nand2 port map( a => n1640, b => n1424, outb => n1639);
   U2198 : xor2 port map( a => n1632, b => n1361, outb => n1637);
   U2199 : oai12 port map( b => n1636, c => n1367, a => n1641, outb => n1632);
   U2200 : aoi22 port map( a => display_out_clk_timer_2_port, b => n1369, c => 
                           display_out_h_row_2_port, d => n1370, outb => n1641)
                           ;
   U2201 : inv port map( inb => display_out_h_col_2_port, outb => n1636);
   U2202 : oai22 port map( a => n1642, b => n1357, c => n424, d => n1358, outb 
                           => display_out_n846);
   U2203 : nand2 port map( a => n1422, b => n1357, outb => n1358);
   U2204 : xor2 port map( a => n1638, b => n1643, outb => n424);
   U2205 : xor2 port map( a => n1361, b => n422, outb => n1643);
   U2206 : inv port map( inb => n1424, outb => n422);
   U2207 : oai12 port map( b => n1423, c => n1367, a => n1644, outb => n1424);
   U2208 : aoi22 port map( a => display_out_clk_timer_0_port, b => n1369, c => 
                           display_out_h_row_0_port, d => n1370, outb => n1644)
                           ;
   U2209 : inv port map( inb => display_out_h_col_0_port, outb => n1423);
   U2210 : inv port map( inb => n1640, outb => n1638);
   U2211 : oai12 port map( b => n1642, c => n1367, a => n1645, outb => n1640);
   U2212 : aoi22 port map( a => display_out_clk_timer_1_port, b => n1369, c => 
                           display_out_h_row_1_port, d => n1370, outb => n1645)
                           ;
   U2213 : inv port map( inb => n1361, outb => n1369);
   U2214 : nor2 port map( a => n1343, b => n1342, outb => n1361);
   U2215 : nand2 port map( a => n1646, b => n1367, outb => n1357);
   U2216 : inv port map( inb => display_out_h_col_1_port, outb => n1642);
   U2217 : oai22 port map( a => n1415, b => n1647, c => n1648, d => n1649, outb
                           => display_out_n845);
   U2218 : inv port map( inb => hub_clk_o_port, outb => n1649);
   U2219 : inv port map( inb => n1648, outb => n1647);
   U2220 : nand2 port map( a => n1650, b => n1418, outb => n1648);
   U2221 : inv port map( inb => n1651, outb => n1418);
   U2222 : nand2 port map( a => n1413, b => n1414, outb => n1651);
   U2223 : aoi12 port map( b => n1652, c => n1343, a => n1653, outb => n1415);
   U2224 : inv port map( inb => n1654, outb => n1653);
   U2225 : nand3 port map( a => n1412, b => n1655, c => n1656, outb => 
                           display_out_n844);
   U2226 : nand3 port map( a => n1411, b => n1421, c => hub_latch_o_port, outb 
                           => n1656);
   U2227 : inv port map( inb => n1657, outb => n1421);
   U2228 : nand2 port map( a => n1345, b => n1342, outb => n1412);
   U2229 : oai22 port map( a => n1658, b => n1659, c => n1660, d => n1655, outb
                           => display_out_n843);
   U2230 : inv port map( inb => n1661, outb => n1660);
   U2231 : oai22 port map( a => n1662, b => n1659, c => 
                           display_out_bcd_time_0_port, d => n1655, outb => 
                           display_out_n842);
   U2232 : inv port map( inb => n1663, outb => n1655);
   U2233 : nand2 port map( a => n1664, b => n1665, outb => display_out_n841);
   U2234 : oai12 port map( b => n1666, c => n1411, a => 
                           display_out_bcd_time_2_port, outb => n1665);
   U2235 : aoi12 port map( b => n1662, c => n1661, a => n1667, outb => n1666);
   U2236 : nand4 port map( a => n1661, b => n1662, c => n1663, d => n1668, outb
                           => n1664);
   U2237 : nor2 port map( a => n1667, b => n1411, outb => n1663);
   U2238 : oai12 port map( b => display_out_bcd_time_1_port, c => 
                           display_out_bcd_time_0_port, a => n1669, outb => 
                           n1661);
   U2239 : nand4 port map( a => n1670, b => n1671, c => n1672, d => n1673, outb
                           => display_out_n840);
   U2240 : nand2 port map( a => n1674, b => n1675, outb => n1671);
   U2241 : aoi22 port map( a => n355, b => n1676, c => n431, d => 
                           display_out_disp_timer_0_port, outb => n1670);
   U2242 : nand3 port map( a => n1677, b => n1678, c => n1679, outb => 
                           display_out_n839);
   U2243 : nand2 port map( a => n355, b => n486, outb => n1679);
   U2244 : oai12 port map( b => display_out_disp_timer_12_port, c => n1680, a 
                           => display_out_disp_timer_13_port, outb => n1677);
   U2245 : nand3 port map( a => n1681, b => n1682, c => n1673, outb => 
                           display_out_n838);
   U2246 : nand2 port map( a => display_out_disp_timer_12_port, b => n1680, 
                           outb => n1682);
   U2247 : nand2 port map( a => n1683, b => n440, outb => n1680);
   U2248 : nand3 port map( a => n355, b => n1683, c => n1684, outb => n1681);
   U2249 : nand3 port map( a => n1685, b => n1686, c => n1687, outb => 
                           display_out_n837);
   U2250 : nand2 port map( a => n355, b => n1683, outb => n1687);
   U2251 : inv port map( inb => n1688, outb => n1683);
   U2252 : inv port map( inb => n1689, outb => n1685);
   U2253 : nor2 port map( a => n1690, b => n1691, outb => n1689);
   U2254 : aoi12 port map( b => n355, c => display_out_disp_timer_10_port, a =>
                           n1692, outb => n1691);
   U2255 : nand3 port map( a => n1693, b => n1694, c => n1695, outb => 
                           display_out_n836);
   U2256 : nand2 port map( a => n1675, b => n1696, outb => n1695);
   U2257 : nand2 port map( a => display_out_disp_timer_10_port, b => n1692, 
                           outb => n1694);
   U2258 : oai12 port map( b => n1697, c => n352, a => n440, outb => n1692);
   U2259 : nand3 port map( a => n355, b => n1697, c => n1698, outb => n1693);
   U2260 : nand3 port map( a => n1699, b => n1678, c => n1700, outb => 
                           display_out_n835);
   U2261 : aoi22 port map( a => n1675, b => n1701, c => n355, d => n1697, outb 
                           => n1700);
   U2262 : oai12 port map( b => display_out_disp_timer_8_port, c => n1702, a =>
                           display_out_disp_timer_9_port, outb => n1699);
   U2263 : nand4 port map( a => n1703, b => n1673, c => n1704, d => n1705, outb
                           => display_out_n834);
   U2264 : nand2 port map( a => display_out_disp_timer_8_port, b => n1702, outb
                           => n1705);
   U2265 : nand2 port map( a => n1706, b => n440, outb => n1702);
   U2266 : nand3 port map( a => n355, b => n1706, c => n1707, outb => n1704);
   U2267 : nand3 port map( a => n1708, b => n1686, c => n1709, outb => 
                           display_out_n833);
   U2268 : aoi22 port map( a => n1675, b => n1710, c => n355, d => n1706, outb 
                           => n1709);
   U2269 : nand2 port map( a => display_out_disp_timer_7_port, b => n1711, outb
                           => n1708);
   U2270 : oai12 port map( b => n1712, c => n352, a => n440, outb => n1711);
   U2271 : nand3 port map( a => n1713, b => n1672, c => n1714, outb => 
                           display_out_n832);
   U2272 : nand2 port map( a => n355, b => n1712, outb => n1714);
   U2273 : nand2 port map( a => display_out_disp_timer_6_port, b => n1715, outb
                           => n1713);
   U2274 : oai12 port map( b => n352, c => n1716, a => n1717, outb => n1715);
   U2275 : nand3 port map( a => n1718, b => n1719, c => n1720, outb => 
                           display_out_n831);
   U2276 : nand2 port map( a => n1675, b => n1701, outb => n1720);
   U2277 : nand2 port map( a => n1721, b => n1722, outb => n1701);
   U2278 : inv port map( inb => n1674, outb => n1721);
   U2279 : nand2 port map( a => display_out_disp_timer_5_port, b => n1723, outb
                           => n1719);
   U2280 : inv port map( inb => n1717, outb => n1723);
   U2281 : aoi12 port map( b => n1724, c => n355, a => n431, outb => n1717);
   U2282 : nand3 port map( a => n355, b => n1725, c => n1716, outb => n1718);
   U2283 : nand4 port map( a => n1726, b => n1727, c => n1678, d => n1703, outb
                           => display_out_n830);
   U2284 : oai12 port map( b => n1674, c => n1728, a => n1675, outb => n1703);
   U2285 : nor3 port map( a => n1662, b => display_out_bcd_time_1_port, c => 
                           n1668, outb => n1674);
   U2286 : nand2 port map( a => n1729, b => n440, outb => n1678);
   U2287 : oai12 port map( b => display_out_disp_timer_3_port, c => n1730, a =>
                           display_out_disp_timer_4_port, outb => n1727);
   U2288 : nand2 port map( a => n355, b => n1725, outb => n1726);
   U2289 : inv port map( inb => n1724, outb => n1725);
   U2290 : nand4 port map( a => n1731, b => n1673, c => n1732, d => n1733, outb
                           => display_out_n829);
   U2291 : nand2 port map( a => display_out_disp_timer_3_port, b => n1730, outb
                           => n1733);
   U2292 : nand2 port map( a => n1734, b => n440, outb => n1730);
   U2293 : nand3 port map( a => n355, b => n1734, c => n1735, outb => n1732);
   U2294 : nand2 port map( a => n1675, b => n1710, outb => n1731);
   U2295 : inv port map( inb => n1736, outb => n1710);
   U2296 : nor2 port map( a => n1737, b => n1728, outb => n1736);
   U2297 : nor3 port map( a => n1658, b => display_out_bcd_time_0_port, c => 
                           n1668, outb => n1728);
   U2298 : nand4 port map( a => n1738, b => n1739, c => n1686, d => n1673, outb
                           => display_out_n828);
   U2299 : nand3 port map( a => display_out_bcd_time_1_port, b => n1668, c => 
                           n1675, outb => n1686);
   U2300 : nor2 port map( a => n1740, b => n431, outb => n1675);
   U2301 : oai12 port map( b => display_out_disp_timer_1_port, c => n1741, a =>
                           display_out_disp_timer_2_port, outb => n1739);
   U2302 : nand2 port map( a => n355, b => n1734, outb => n1738);
   U2303 : nand4 port map( a => n1672, b => n1673, c => n1742, d => n1743, outb
                           => display_out_n827);
   U2304 : nand2 port map( a => display_out_disp_timer_1_port, b => n1741, outb
                           => n1743);
   U2305 : nand2 port map( a => n440, b => n1676, outb => n1741);
   U2306 : nand3 port map( a => n355, b => n1676, c => n1744, outb => n1742);
   U2307 : inv port map( inb => n352, outb => n355);
   U2308 : oai12 port map( b => n1745, c => n1374, a => n440, outb => n352);
   U2309 : nand2 port map( a => n1746, b => n1747, outb => n1374);
   U2310 : inv port map( inb => n1339, outb => n1745);
   U2311 : nand2 port map( a => n1748, b => n440, outb => n1673);
   U2312 : nand2 port map( a => n1749, b => n1750, outb => n1748);
   U2313 : nand4 port map( a => display_out_bcd_time_1_port, b => n1350, c => 
                           n1662, d => n1668, outb => n1750);
   U2314 : inv port map( inb => n1729, outb => n1749);
   U2315 : nand2 port map( a => n1646, b => n1751, outb => n1729);
   U2316 : nand4 port map( a => display_out_bcd_time_0_port, b => n1350, c => 
                           n1658, d => n1668, outb => n1751);
   U2317 : inv port map( inb => n1752, outb => n1672);
   U2318 : nor3 port map( a => n1753, b => n431, c => n1740, outb => n1752);
   U2319 : inv port map( inb => n440, outb => n431);
   U2320 : nand4 port map( a => n1419, b => n1746, c => n1413, d => n1646, outb
                           => n440);
   U2321 : oai12 port map( b => n1342, c => n1754, a => n1422, outb => n1413);
   U2322 : inv port map( inb => n1755, outb => n1754);
   U2323 : inv port map( inb => n1756, outb => n1419);
   U2324 : oai12 port map( b => n1667, c => n351, a => n1339, outb => n1756);
   U2325 : nand2 port map( a => n1342, b => n1404, outb => n1339);
   U2326 : nor2 port map( a => n1696, b => n1737, outb => n1753);
   U2327 : oai12 port map( b => display_out_bcd_time_2_port, c => n1669, a => 
                           n1722, outb => n1696);
   U2328 : nand3 port map( a => n1662, b => n1658, c => 
                           display_out_bcd_time_2_port, outb => n1722);
   U2329 : inv port map( inb => display_out_bcd_time_1_port, outb => n1658);
   U2330 : inv port map( inb => display_out_bcd_time_0_port, outb => n1662);
   U2331 : oai12 port map( b => n1650, c => n1757, a => n1758, outb => 
                           display_out_n826);
   U2332 : nand2 port map( a => hub_blank_o_port, b => n1757, outb => n1758);
   U2333 : nor2 port map( a => n358, b => n1657, outb => n1757);
   U2334 : inv port map( inb => n416, outb => n358);
   U2335 : nand3 port map( a => n1759, b => n1646, c => n1760, outb => 
                           display_out_n825);
   U2336 : nand2 port map( a => hub_mux_o_0_port, b => n416, outb => n1760);
   U2337 : nand2 port map( a => n418, b => display_out_h_row_0_port, outb => 
                           n1759);
   U2338 : nand3 port map( a => n1761, b => n1646, c => n1762, outb => 
                           display_out_n824);
   U2339 : nand2 port map( a => hub_mux_o_1_port, b => n416, outb => n1762);
   U2340 : nand2 port map( a => n418, b => display_out_h_row_1_port, outb => 
                           n1761);
   U2341 : nand3 port map( a => n1763, b => n1646, c => n1764, outb => 
                           display_out_n823);
   U2342 : nand2 port map( a => hub_mux_o_2_port, b => n416, outb => n1764);
   U2343 : nand2 port map( a => n418, b => display_out_h_row_2_port, outb => 
                           n1763);
   U2344 : nand3 port map( a => n1765, b => n1646, c => n1766, outb => 
                           display_out_n822);
   U2345 : nand2 port map( a => hub_mux_o_3_port, b => n416, outb => n1766);
   U2346 : nand2 port map( a => n418, b => display_out_h_row_3_port, outb => 
                           n1765);
   U2347 : nor2 port map( a => n1667, b => n416, outb => n418);
   U2348 : nor2 port map( a => n1370, b => n1346, outb => n416);
   U2349 : inv port map( inb => n1767, outb => n1370);
   U2350 : nand2 port map( a => n1768, b => n1737, outb => n1767);
   U2351 : nor2 port map( a => n1668, b => n1669, outb => n1737);
   U2352 : nand2 port map( a => display_out_bcd_time_1_port, b => 
                           display_out_bcd_time_0_port, outb => n1669);
   U2353 : inv port map( inb => display_out_bcd_time_2_port, outb => n1668);
   U2354 : oai22 port map( a => n1769, b => n1770, c => n56, d => n1771, outb 
                           => display_out_n821);
   U2355 : inv port map( inb => hub_reg_f, outb => n56);
   U2356 : aoi12 port map( b => n1344, c => n1346, a => n1345, outb => n1770);
   U2357 : inv port map( inb => n1771, outb => n1769);
   U2358 : nand3 port map( a => n1772, b => n1646, c => n1773, outb => n1771);
   U2359 : nand2 port map( a => n1657, b => n1344, outb => n1773);
   U2360 : nor2 port map( a => n1352, b => n1755, outb => n1657);
   U2361 : inv port map( inb => n1345, outb => n1352);
   U2362 : inv port map( inb => n1346, outb => n1646);
   U2363 : nand2 port map( a => n1342, b => n1343, outb => n1772);
   U2364 : oai12 port map( b => n1774, c => n1775, a => n1776, outb => 
                           display_out_n820);
   U2365 : aoi22 port map( a => display_out_hub_piso_r0_2_port, b => n1777, c 
                           => n1778, d => mem_sipo_r0_1_port, outb => n1776);
   U2366 : inv port map( inb => display_out_hub_piso_r0_1_port, outb => n1775);
   U2367 : oai12 port map( b => n1779, c => n1774, a => n1780, outb => 
                           display_out_n819);
   U2368 : aoi22 port map( a => display_out_hub_piso_r0_3_port, b => n1777, c 
                           => n1778, d => mem_sipo_r0_2_port, outb => n1780);
   U2369 : inv port map( inb => display_out_hub_piso_r0_2_port, outb => n1779);
   U2370 : oai12 port map( b => n1774, c => n1781, a => n1782, outb => 
                           display_out_n818);
   U2371 : aoi22 port map( a => display_out_hub_piso_r0_4_port, b => n1777, c 
                           => n1778, d => mem_sipo_r0_3_port, outb => n1782);
   U2372 : inv port map( inb => display_out_hub_piso_r0_3_port, outb => n1781);
   U2373 : oai12 port map( b => n1774, c => n1783, a => n1784, outb => 
                           display_out_n817);
   U2374 : aoi22 port map( a => display_out_hub_piso_r0_5_port, b => n1777, c 
                           => n1778, d => mem_sipo_r0_4_port, outb => n1784);
   U2375 : inv port map( inb => display_out_hub_piso_r0_4_port, outb => n1783);
   U2376 : oai12 port map( b => n1774, c => n1785, a => n1786, outb => 
                           display_out_n816);
   U2377 : aoi22 port map( a => display_out_hub_piso_r0_6_port, b => n1777, c 
                           => n1778, d => mem_sipo_r0_5_port, outb => n1786);
   U2378 : inv port map( inb => display_out_hub_piso_r0_5_port, outb => n1785);
   U2379 : oai12 port map( b => n1774, c => n1787, a => n1788, outb => 
                           display_out_n815);
   U2380 : aoi22 port map( a => n1777, b => display_out_hub_piso_r0_7_port, c 
                           => n1778, d => mem_sipo_r0_6_port, outb => n1788);
   U2381 : inv port map( inb => display_out_hub_piso_r0_6_port, outb => n1787);
   U2382 : oai12 port map( b => n1774, c => n1789, a => n1790, outb => 
                           display_out_n814);
   U2383 : aoi22 port map( a => display_out_hub_piso_r0_1_port, b => n1777, c 
                           => n1778, d => mem_sipo_r0_0_port, outb => n1790);
   U2384 : oai12 port map( b => n1774, c => n1791, a => n1792, outb => 
                           display_out_n813);
   U2385 : aoi22 port map( a => display_out_hub_piso_g0_2_port, b => n1777, c 
                           => n1778, d => mem_sipo_g0_1_port, outb => n1792);
   U2386 : inv port map( inb => display_out_hub_piso_g0_1_port, outb => n1791);
   U2387 : oai12 port map( b => n1774, c => n1793, a => n1794, outb => 
                           display_out_n812);
   U2388 : aoi22 port map( a => display_out_hub_piso_g0_3_port, b => n1777, c 
                           => n1778, d => mem_sipo_g0_2_port, outb => n1794);
   U2389 : inv port map( inb => display_out_hub_piso_g0_2_port, outb => n1793);
   U2390 : oai12 port map( b => n1774, c => n1795, a => n1796, outb => 
                           display_out_n811);
   U2391 : aoi22 port map( a => display_out_hub_piso_g0_4_port, b => n1777, c 
                           => n1778, d => mem_sipo_g0_3_port, outb => n1796);
   U2392 : inv port map( inb => display_out_hub_piso_g0_3_port, outb => n1795);
   U2393 : oai12 port map( b => n1774, c => n1797, a => n1798, outb => 
                           display_out_n810);
   U2394 : aoi22 port map( a => display_out_hub_piso_g0_5_port, b => n1777, c 
                           => n1778, d => mem_sipo_g0_4_port, outb => n1798);
   U2395 : inv port map( inb => display_out_hub_piso_g0_4_port, outb => n1797);
   U2396 : oai12 port map( b => n1774, c => n1799, a => n1800, outb => 
                           display_out_n809);
   U2397 : aoi22 port map( a => display_out_hub_piso_g0_6_port, b => n1777, c 
                           => n1778, d => mem_sipo_g0_5_port, outb => n1800);
   U2398 : inv port map( inb => display_out_hub_piso_g0_5_port, outb => n1799);
   U2399 : oai12 port map( b => n1774, c => n1801, a => n1802, outb => 
                           display_out_n808);
   U2400 : aoi22 port map( a => n1777, b => display_out_hub_piso_g0_7_port, c 
                           => n1778, d => mem_sipo_g0_6_port, outb => n1802);
   U2401 : inv port map( inb => display_out_hub_piso_g0_6_port, outb => n1801);
   U2402 : oai12 port map( b => n1774, c => n1803, a => n1804, outb => 
                           display_out_n807);
   U2403 : aoi22 port map( a => display_out_hub_piso_g0_1_port, b => n1777, c 
                           => n1778, d => mem_sipo_g0_0_port, outb => n1804);
   U2404 : oai12 port map( b => n1774, c => n1805, a => n1806, outb => 
                           display_out_n806);
   U2405 : aoi22 port map( a => display_out_hub_piso_b0_2_port, b => n1777, c 
                           => n1778, d => mem_sipo_b0_1_port, outb => n1806);
   U2406 : inv port map( inb => display_out_hub_piso_b0_1_port, outb => n1805);
   U2407 : oai12 port map( b => n1774, c => n1807, a => n1808, outb => 
                           display_out_n805);
   U2408 : aoi22 port map( a => display_out_hub_piso_b0_3_port, b => n1777, c 
                           => n1778, d => mem_sipo_b0_2_port, outb => n1808);
   U2409 : inv port map( inb => display_out_hub_piso_b0_2_port, outb => n1807);
   U2410 : oai12 port map( b => n1774, c => n1809, a => n1810, outb => 
                           display_out_n804);
   U2411 : aoi22 port map( a => display_out_hub_piso_b0_4_port, b => n1777, c 
                           => n1778, d => mem_sipo_b0_3_port, outb => n1810);
   U2412 : inv port map( inb => display_out_hub_piso_b0_3_port, outb => n1809);
   U2413 : oai12 port map( b => n1774, c => n1811, a => n1812, outb => 
                           display_out_n803);
   U2414 : aoi22 port map( a => display_out_hub_piso_b0_5_port, b => n1777, c 
                           => n1778, d => mem_sipo_b0_4_port, outb => n1812);
   U2415 : inv port map( inb => display_out_hub_piso_b0_4_port, outb => n1811);
   U2416 : oai12 port map( b => n1774, c => n1813, a => n1814, outb => 
                           display_out_n802);
   U2417 : aoi22 port map( a => display_out_hub_piso_b0_6_port, b => n1777, c 
                           => n1778, d => mem_sipo_b0_5_port, outb => n1814);
   U2418 : inv port map( inb => display_out_hub_piso_b0_5_port, outb => n1813);
   U2419 : oai12 port map( b => n1774, c => n1815, a => n1816, outb => 
                           display_out_n801);
   U2420 : aoi22 port map( a => n1777, b => display_out_hub_piso_b0_7_port, c 
                           => n1778, d => mem_sipo_b0_6_port, outb => n1816);
   U2421 : inv port map( inb => display_out_hub_piso_b0_6_port, outb => n1815);
   U2422 : oai12 port map( b => n1774, c => n1817, a => n1818, outb => 
                           display_out_n800);
   U2423 : aoi22 port map( a => display_out_hub_piso_b0_1_port, b => n1777, c 
                           => n1778, d => mem_sipo_b0_0_port, outb => n1818);
   U2424 : nor2 port map( a => n1650, b => n1819, outb => n1778);
   U2425 : nor2 port map( a => n1346, b => n1404, outb => n1650);
   U2426 : nor2 port map( a => n1747, b => n1819, outb => n1777);
   U2427 : inv port map( inb => n1774, outb => n1819);
   U2428 : nand2 port map( a => n1367, b => n339, outb => n1774);
   U2429 : oai12 port map( b => n1768, c => n1344, a => n1659, outb => n339);
   U2430 : inv port map( inb => n1411, outb => n1659);
   U2431 : nor2 port map( a => n1346, b => n1768, outb => n1411);
   U2432 : nor3 port map( a => display_out_hub_out_sm_1_port, b => 
                           display_out_hub_out_sm_2_port, c => 
                           display_out_hub_out_sm_0_port, outb => n1346);
   U2433 : nor2 port map( a => n501, b => n1820, outb => n1344);
   U2434 : inv port map( inb => reg_hub_f, outb => n1820);
   U2435 : inv port map( inb => mem_hub_f, outb => n501);
   U2436 : nor2 port map( a => n351, b => n1740, outb => n1768);
   U2437 : inv port map( inb => n1350, outb => n1740);
   U2438 : nor2 port map( a => n1667, b => n1342, outb => n1350);
   U2439 : inv port map( inb => n1652, outb => n1342);
   U2440 : nand4 port map( a => n434, b => n428, c => n1821, d => n354, outb =>
                           n351);
   U2441 : inv port map( inb => display_out_disp_timer_31_port, outb => n354);
   U2442 : inv port map( inb => display_out_disp_timer_30_port, outb => n1821);
   U2443 : inv port map( inb => display_out_disp_timer_29_port, outb => n428);
   U2444 : inv port map( inb => n430, outb => n434);
   U2445 : nand3 port map( a => n437, b => n433, c => n439, outb => n430);
   U2446 : nor3 port map( a => display_out_disp_timer_25_port, b => 
                           display_out_disp_timer_26_port, c => n447, outb => 
                           n439);
   U2447 : nand2 port map( a => n451, b => n450, outb => n447);
   U2448 : inv port map( inb => display_out_disp_timer_24_port, outb => n450);
   U2449 : nor3 port map( a => display_out_disp_timer_22_port, b => 
                           display_out_disp_timer_23_port, c => n458, outb => 
                           n451);
   U2450 : nand3 port map( a => n463, b => n460, c => n465, outb => n458);
   U2451 : nor3 port map( a => display_out_disp_timer_18_port, b => 
                           display_out_disp_timer_19_port, c => n472, outb => 
                           n465);
   U2452 : inv port map( inb => n471, outb => n472);
   U2453 : nor3 port map( a => display_out_disp_timer_16_port, b => 
                           display_out_disp_timer_17_port, c => n479, outb => 
                           n471);
   U2454 : nand3 port map( a => n484, b => n481, c => n486, outb => n479);
   U2455 : nor3 port map( a => display_out_disp_timer_12_port, b => 
                           display_out_disp_timer_13_port, c => n1688, outb => 
                           n486);
   U2456 : nand3 port map( a => n1698, b => n1690, c => n1697, outb => n1688);
   U2457 : nor3 port map( a => display_out_disp_timer_8_port, b => 
                           display_out_disp_timer_9_port, c => n1822, outb => 
                           n1697);
   U2458 : inv port map( inb => n1706, outb => n1822);
   U2459 : nor2 port map( a => n1823, b => display_out_disp_timer_7_port, outb 
                           => n1706);
   U2460 : inv port map( inb => n1712, outb => n1823);
   U2461 : nor3 port map( a => display_out_disp_timer_5_port, b => 
                           display_out_disp_timer_6_port, c => n1724, outb => 
                           n1712);
   U2462 : nand3 port map( a => n1735, b => n1824, c => n1734, outb => n1724);
   U2463 : nor3 port map( a => display_out_disp_timer_1_port, b => 
                           display_out_disp_timer_2_port, c => 
                           display_out_disp_timer_0_port, outb => n1734);
   U2464 : nand2 port map( a => n1406, b => n1652, outb => n1367);
   U2465 : nand3 port map( a => n1825, b => n1826, c => n1827, outb => n1652);
   U2466 : aoi22 port map( a => display_out_h_col_31_port, b => n1406, c => 
                           display_out_clk_timer_31_port, d => n1410, outb => 
                           n1827);
   U2467 : nand2 port map( a => display_out_disp_timer_31_port, b => n1404, 
                           outb => n1826);
   U2468 : nand4 port map( a => n1828, b => n1829, c => n1830, d => n1831, outb
                           => n1825);
   U2469 : aoi22 port map( a => n1406, b => n1832, c => n1833, d => n1414, outb
                           => n1831);
   U2470 : nand4 port map( a => n1834, b => n1835, c => n1836, d => n1837, outb
                           => n1832);
   U2471 : nor2 port map( a => n1838, b => n1839, outb => n1837);
   U2472 : nand3 port map( a => n1621, b => n1613, c => n1629, outb => n1839);
   U2473 : inv port map( inb => display_out_h_col_3_port, outb => n1629);
   U2474 : inv port map( inb => display_out_h_col_5_port, outb => n1613);
   U2475 : inv port map( inb => display_out_h_col_4_port, outb => n1621);
   U2476 : nand4 port map( a => n1606, b => n1599, c => n1590, d => n1583, outb
                           => n1838);
   U2477 : inv port map( inb => display_out_h_col_9_port, outb => n1583);
   U2478 : inv port map( inb => display_out_h_col_8_port, outb => n1590);
   U2479 : inv port map( inb => display_out_h_col_7_port, outb => n1599);
   U2480 : inv port map( inb => display_out_h_col_6_port, outb => n1606);
   U2481 : nor2 port map( a => n1840, b => n1841, outb => n1836);
   U2482 : nand3 port map( a => n1463, b => n1455, c => n1471, outb => n1841);
   U2483 : inv port map( inb => display_out_h_col_24_port, outb => n1471);
   U2484 : inv port map( inb => display_out_h_col_26_port, outb => n1455);
   U2485 : inv port map( inb => display_out_h_col_25_port, outb => n1463);
   U2486 : nand4 port map( a => n1448, b => n1440, c => n1433, d => n1425, outb
                           => n1840);
   U2487 : inv port map( inb => display_out_h_col_30_port, outb => n1425);
   U2488 : inv port map( inb => display_out_h_col_29_port, outb => n1433);
   U2489 : inv port map( inb => display_out_h_col_28_port, outb => n1440);
   U2490 : inv port map( inb => display_out_h_col_27_port, outb => n1448);
   U2491 : nor2 port map( a => n1842, b => n1843, outb => n1835);
   U2492 : nand3 port map( a => n1516, b => n1508, c => n1523, outb => n1843);
   U2493 : inv port map( inb => display_out_h_col_17_port, outb => n1523);
   U2494 : inv port map( inb => display_out_h_col_19_port, outb => n1508);
   U2495 : inv port map( inb => display_out_h_col_18_port, outb => n1516);
   U2496 : nand4 port map( a => n1501, b => n1493, c => n1486, d => n1478, outb
                           => n1842);
   U2497 : inv port map( inb => display_out_h_col_23_port, outb => n1478);
   U2498 : inv port map( inb => display_out_h_col_22_port, outb => n1486);
   U2499 : inv port map( inb => display_out_h_col_21_port, outb => n1493);
   U2500 : inv port map( inb => display_out_h_col_20_port, outb => n1501);
   U2501 : nor2 port map( a => n1844, b => n1845, outb => n1834);
   U2502 : nand3 port map( a => n1568, b => n1561, c => n1575, outb => n1845);
   U2503 : inv port map( inb => display_out_h_col_10_port, outb => n1575);
   U2504 : inv port map( inb => display_out_h_col_12_port, outb => n1561);
   U2505 : inv port map( inb => display_out_h_col_11_port, outb => n1568);
   U2506 : nand4 port map( a => n1553, b => n1546, c => n1538, d => n1531, outb
                           => n1844);
   U2507 : inv port map( inb => display_out_h_col_16_port, outb => n1531);
   U2508 : inv port map( inb => display_out_h_col_15_port, outb => n1538);
   U2509 : inv port map( inb => display_out_h_col_14_port, outb => n1546);
   U2510 : inv port map( inb => display_out_h_col_13_port, outb => n1553);
   U2511 : oai12 port map( b => n1846, c => n1847, a => n1410, outb => n1830);
   U2512 : oai12 port map( b => n1833, c => n1414, a => n1848, outb => n1829);
   U2513 : inv port map( inb => n1849, outb => n1848);
   U2514 : oai22 port map( a => n1338, b => n1850, c => n1851, d => n1852, outb
                           => n1849);
   U2515 : inv port map( inb => n1853, outb => n1850);
   U2516 : nand2 port map( a => n1851, b => n1852, outb => n1853);
   U2517 : oai12 port map( b => n1667, c => n1676, a => n1854, outb => n1852);
   U2518 : aoi22 port map( a => display_out_h_col_0_port, b => n1406, c => 
                           display_out_clk_timer_0_port, d => n1410, outb => 
                           n1854);
   U2519 : inv port map( inb => display_out_disp_timer_0_port, outb => n1676);
   U2520 : oai12 port map( b => n1667, c => n1744, a => n1855, outb => n1851);
   U2521 : aoi22 port map( a => display_out_h_col_1_port, b => n1406, c => 
                           display_out_clk_timer_1_port, d => n1410, outb => 
                           n1855);
   U2522 : inv port map( inb => display_out_disp_timer_1_port, outb => n1744);
   U2523 : inv port map( inb => n1406, outb => n1338);
   U2524 : oai12 port map( b => n1667, c => n1856, a => n1857, outb => n1833);
   U2525 : aoi22 port map( a => display_out_h_col_2_port, b => n1406, c => 
                           display_out_clk_timer_2_port, d => n1410, outb => 
                           n1857);
   U2526 : nand2 port map( a => n1746, b => n1654, outb => n1410);
   U2527 : nand2 port map( a => n1422, b => n1755, outb => n1654);
   U2528 : inv port map( inb => n1747, outb => n1422);
   U2529 : nor2 port map( a => n1343, b => n1345, outb => n1746);
   U2530 : nor3 port map( a => display_out_hub_out_sm_0_port, b => 
                           display_out_hub_out_sm_1_port, c => n1349, outb => 
                           n1345);
   U2531 : inv port map( inb => display_out_disp_timer_2_port, outb => n1856);
   U2532 : nand2 port map( a => n1404, b => n1858, outb => n1828);
   U2533 : nand2 port map( a => n1859, b => n1860, outb => n1858);
   U2534 : nor3 port map( a => n1861, b => n1862, c => n1863, outb => n1860);
   U2535 : nand3 port map( a => n1824, b => n1716, c => n1735, outb => n1863);
   U2536 : inv port map( inb => display_out_disp_timer_3_port, outb => n1735);
   U2537 : inv port map( inb => display_out_disp_timer_5_port, outb => n1716);
   U2538 : inv port map( inb => display_out_disp_timer_4_port, outb => n1824);
   U2539 : nand4 port map( a => n1864, b => n1865, c => n1707, d => n1866, outb
                           => n1862);
   U2540 : inv port map( inb => display_out_disp_timer_9_port, outb => n1866);
   U2541 : inv port map( inb => display_out_disp_timer_8_port, outb => n1707);
   U2542 : inv port map( inb => display_out_disp_timer_7_port, outb => n1865);
   U2543 : inv port map( inb => display_out_disp_timer_6_port, outb => n1864);
   U2544 : nand4 port map( a => n437, b => n433, c => n1867, d => n1868, outb 
                           => n1861);
   U2545 : nor3 port map( a => display_out_disp_timer_24_port, b => 
                           display_out_disp_timer_26_port, c => 
                           display_out_disp_timer_25_port, outb => n1868);
   U2546 : nor2 port map( a => display_out_disp_timer_30_port, b => 
                           display_out_disp_timer_29_port, outb => n1867);
   U2547 : inv port map( inb => display_out_disp_timer_28_port, outb => n433);
   U2548 : inv port map( inb => display_out_disp_timer_27_port, outb => n437);
   U2549 : nor3 port map( a => n1869, b => n1870, c => n1871, outb => n1859);
   U2550 : nand3 port map( a => n1690, b => n1684, c => n1698, outb => n1871);
   U2551 : inv port map( inb => display_out_disp_timer_10_port, outb => n1698);
   U2552 : inv port map( inb => display_out_disp_timer_12_port, outb => n1684);
   U2553 : inv port map( inb => display_out_disp_timer_11_port, outb => n1690);
   U2554 : nand4 port map( a => n1872, b => n484, c => n481, d => n475, outb =>
                           n1870);
   U2555 : inv port map( inb => display_out_disp_timer_16_port, outb => n475);
   U2556 : inv port map( inb => display_out_disp_timer_15_port, outb => n481);
   U2557 : inv port map( inb => display_out_disp_timer_14_port, outb => n484);
   U2558 : inv port map( inb => display_out_disp_timer_13_port, outb => n1872);
   U2559 : nand4 port map( a => n463, b => n460, c => n1873, d => n1874, outb 
                           => n1869);
   U2560 : nor3 port map( a => display_out_disp_timer_17_port, b => 
                           display_out_disp_timer_19_port, c => 
                           display_out_disp_timer_18_port, outb => n1874);
   U2561 : nor2 port map( a => display_out_disp_timer_23_port, b => 
                           display_out_disp_timer_22_port, outb => n1873);
   U2562 : inv port map( inb => display_out_disp_timer_21_port, outb => n460);
   U2563 : inv port map( inb => display_out_disp_timer_20_port, outb => n463);
   U2564 : inv port map( inb => n1667, outb => n1404);
   U2565 : nand3 port map( a => display_out_hub_out_sm_1_port, b => n1349, c =>
                           display_out_hub_out_sm_0_port, outb => n1667);
   U2566 : nor2 port map( a => n1747, b => n1755, outb => n1406);
   U2567 : nand4 port map( a => n1875, b => n1373, c => n1876, d => n1877, outb
                           => n1755);
   U2568 : nor3 port map( a => display_out_clk_timer_1_port, b => 
                           display_out_clk_timer_31_port, c => 
                           display_out_clk_timer_2_port, outb => n1877);
   U2569 : inv port map( inb => n1847, outb => n1876);
   U2570 : nand3 port map( a => n1878, b => n1879, c => n1880, outb => n1847);
   U2571 : nor2 port map( a => n1881, b => n1882, outb => n1880);
   U2572 : nand3 port map( a => n1390, b => n1389, c => n1391, outb => n1882);
   U2573 : inv port map( inb => display_out_clk_timer_16_port, outb => n1391);
   U2574 : inv port map( inb => display_out_clk_timer_18_port, outb => n1389);
   U2575 : inv port map( inb => display_out_clk_timer_17_port, outb => n1390);
   U2576 : nand4 port map( a => n1388, b => n1387, c => n1386, d => n1385, outb
                           => n1881);
   U2577 : inv port map( inb => display_out_clk_timer_22_port, outb => n1385);
   U2578 : inv port map( inb => display_out_clk_timer_21_port, outb => n1386);
   U2579 : inv port map( inb => display_out_clk_timer_20_port, outb => n1387);
   U2580 : inv port map( inb => display_out_clk_timer_19_port, outb => n1388);
   U2581 : nor3 port map( a => display_out_clk_timer_13_port, b => 
                           display_out_clk_timer_15_port, c => 
                           display_out_clk_timer_14_port, outb => n1879);
   U2582 : nor3 port map( a => display_out_clk_timer_10_port, b => 
                           display_out_clk_timer_12_port, c => 
                           display_out_clk_timer_11_port, outb => n1878);
   U2583 : inv port map( inb => display_out_clk_timer_0_port, outb => n1373);
   U2584 : inv port map( inb => n1846, outb => n1875);
   U2585 : nand2 port map( a => n1883, b => n1884, outb => n1846);
   U2586 : nor2 port map( a => n1885, b => n1886, outb => n1884);
   U2587 : nand4 port map( a => n1377, b => n1887, c => n1888, d => n1402, outb
                           => n1886);
   U2588 : inv port map( inb => display_out_clk_timer_5_port, outb => n1402);
   U2589 : inv port map( inb => display_out_clk_timer_4_port, outb => n1888);
   U2590 : inv port map( inb => display_out_clk_timer_3_port, outb => n1887);
   U2591 : inv port map( inb => display_out_clk_timer_30_port, outb => n1377);
   U2592 : nand4 port map( a => n1401, b => n1400, c => n1399, d => n1398, outb
                           => n1885);
   U2593 : inv port map( inb => display_out_clk_timer_9_port, outb => n1398);
   U2594 : inv port map( inb => display_out_clk_timer_8_port, outb => n1399);
   U2595 : inv port map( inb => display_out_clk_timer_7_port, outb => n1400);
   U2596 : inv port map( inb => display_out_clk_timer_6_port, outb => n1401);
   U2597 : nor2 port map( a => n1889, b => n1890, outb => n1883);
   U2598 : nand3 port map( a => n1383, b => n1382, c => n1384, outb => n1890);
   U2599 : inv port map( inb => display_out_clk_timer_23_port, outb => n1384);
   U2600 : inv port map( inb => display_out_clk_timer_25_port, outb => n1382);
   U2601 : inv port map( inb => display_out_clk_timer_24_port, outb => n1383);
   U2602 : nand4 port map( a => n1381, b => n1380, c => n1379, d => n1378, outb
                           => n1889);
   U2603 : inv port map( inb => display_out_clk_timer_29_port, outb => n1378);
   U2604 : inv port map( inb => display_out_clk_timer_28_port, outb => n1379);
   U2605 : inv port map( inb => display_out_clk_timer_27_port, outb => n1380);
   U2606 : inv port map( inb => display_out_clk_timer_26_port, outb => n1381);
   U2607 : nand3 port map( a => n1334, b => n1349, c => 
                           display_out_hub_out_sm_1_port, outb => n1747);
   U2608 : inv port map( inb => display_out_hub_out_sm_2_port, outb => n1349);
   U2609 : oai12 port map( b => n1414, c => n1789, a => n1891, outb => 
                           display_out_n799);
   U2610 : nand2 port map( a => hub_r0_o_port, b => n1414, outb => n1891);
   U2611 : inv port map( inb => display_out_hub_piso_r0_0_port, outb => n1789);
   U2612 : oai12 port map( b => n1414, c => n1803, a => n1892, outb => 
                           display_out_n798);
   U2613 : nand2 port map( a => hub_g0_o_port, b => n1414, outb => n1892);
   U2614 : inv port map( inb => display_out_hub_piso_g0_0_port, outb => n1803);
   U2615 : oai12 port map( b => n1414, c => n1817, a => n1893, outb => 
                           display_out_n797);
   U2616 : nand2 port map( a => hub_b0_o_port, b => n1414, outb => n1893);
   U2617 : inv port map( inb => display_out_hub_piso_b0_0_port, outb => n1817);
   U2618 : inv port map( inb => n1343, outb => n1414);
   U2619 : nor3 port map( a => display_out_hub_out_sm_1_port, b => 
                           display_out_hub_out_sm_2_port, c => n1334, outb => 
                           n1343);
   U2620 : inv port map( inb => display_out_hub_out_sm_0_port, outb => n1334);

end SYN_rtl;
